//
// Verilog description for cell ordenador, 
// 06/12/24 10:25:41
//
// LeonardoSpectrum Level 3, 2020a.2 
//


module ordenador ( y8, y7, y6, y5, y4, y3, y2, y1, x8, x7, x6, x5, x4, x3, x2, 
                   x1 ) ;

    output [63:0]y8 ;
    output [63:0]y7 ;
    output [63:0]y6 ;
    output [63:0]y5 ;
    output [63:0]y4 ;
    output [63:0]y3 ;
    output [63:0]y2 ;
    output [63:0]y1 ;
    input [63:0]x8 ;
    input [63:0]x7 ;
    input [63:0]x6 ;
    input [63:0]x5 ;
    input [63:0]x4 ;
    input [63:0]x3 ;
    input [63:0]x2 ;
    input [63:0]x1 ;

    wire linha7_7__63, linha7_7__62, linha7_7__61, linha7_7__60, linha7_7__59, 
         linha7_7__58, linha7_7__57, linha7_7__56, linha7_7__55, linha7_7__54, 
         linha7_7__53, linha7_7__52, linha7_7__51, linha7_7__50, linha7_7__49, 
         linha7_7__48, linha7_7__47, linha7_7__46, linha7_7__45, linha7_7__44, 
         linha7_7__43, linha7_7__42, linha7_7__41, linha7_7__40, linha7_7__39, 
         linha7_7__38, linha7_7__37, linha7_7__36, linha7_7__35, linha7_7__34, 
         linha7_7__33, linha7_7__32, linha7_7__31, linha7_7__30, linha7_7__29, 
         linha7_7__28, linha7_7__27, linha7_7__26, linha7_7__25, linha7_7__24, 
         linha7_7__23, linha7_7__22, linha7_7__21, linha7_7__20, linha7_7__19, 
         linha7_7__18, linha7_7__17, linha7_7__16, linha7_7__15, linha7_7__14, 
         linha7_7__13, linha7_7__12, linha7_7__11, linha7_7__10, linha7_7__9, 
         linha7_7__8, linha7_7__7, linha7_7__6, linha7_7__5, linha7_7__4, 
         linha7_7__3, linha7_7__2, linha7_7__1, linha7_7__0, linha7_6__63, 
         linha7_6__62, linha7_6__61, linha7_6__60, linha7_6__59, linha7_6__58, 
         linha7_6__57, linha7_6__56, linha7_6__55, linha7_6__54, linha7_6__53, 
         linha7_6__52, linha7_6__51, linha7_6__50, linha7_6__49, linha7_6__48, 
         linha7_6__47, linha7_6__46, linha7_6__45, linha7_6__44, linha7_6__43, 
         linha7_6__42, linha7_6__41, linha7_6__40, linha7_6__39, linha7_6__38, 
         linha7_6__37, linha7_6__36, linha7_6__35, linha7_6__34, linha7_6__33, 
         linha7_6__32, linha7_6__31, linha7_6__30, linha7_6__29, linha7_6__28, 
         linha7_6__27, linha7_6__26, linha7_6__25, linha7_6__24, linha7_6__23, 
         linha7_6__22, linha7_6__21, linha7_6__20, linha7_6__19, linha7_6__18, 
         linha7_6__17, linha7_6__16, linha7_6__15, linha7_6__14, linha7_6__13, 
         linha7_6__12, linha7_6__11, linha7_6__10, linha7_6__9, linha7_6__8, 
         linha7_6__7, linha7_6__6, linha7_6__5, linha7_6__4, linha7_6__3, 
         linha7_6__2, linha7_6__1, linha7_6__0, linha7_5__63, linha7_5__62, 
         linha7_5__61, linha7_5__60, linha7_5__59, linha7_5__58, linha7_5__57, 
         linha7_5__56, linha7_5__55, linha7_5__54, linha7_5__53, linha7_5__52, 
         linha7_5__51, linha7_5__50, linha7_5__49, linha7_5__48, linha7_5__47, 
         linha7_5__46, linha7_5__45, linha7_5__44, linha7_5__43, linha7_5__42, 
         linha7_5__41, linha7_5__40, linha7_5__39, linha7_5__38, linha7_5__37, 
         linha7_5__36, linha7_5__35, linha7_5__34, linha7_5__33, linha7_5__32, 
         linha7_5__31, linha7_5__30, linha7_5__29, linha7_5__28, linha7_5__27, 
         linha7_5__26, linha7_5__25, linha7_5__24, linha7_5__23, linha7_5__22, 
         linha7_5__21, linha7_5__20, linha7_5__19, linha7_5__18, linha7_5__17, 
         linha7_5__16, linha7_5__15, linha7_5__14, linha7_5__13, linha7_5__12, 
         linha7_5__11, linha7_5__10, linha7_5__9, linha7_5__8, linha7_5__7, 
         linha7_5__6, linha7_5__5, linha7_5__4, linha7_5__3, linha7_5__2, 
         linha7_5__1, linha7_5__0, linha7_4__63, linha7_4__62, linha7_4__61, 
         linha7_4__60, linha7_4__59, linha7_4__58, linha7_4__57, linha7_4__56, 
         linha7_4__55, linha7_4__54, linha7_4__53, linha7_4__52, linha7_4__51, 
         linha7_4__50, linha7_4__49, linha7_4__48, linha7_4__47, linha7_4__46, 
         linha7_4__45, linha7_4__44, linha7_4__43, linha7_4__42, linha7_4__41, 
         linha7_4__40, linha7_4__39, linha7_4__38, linha7_4__37, linha7_4__36, 
         linha7_4__35, linha7_4__34, linha7_4__33, linha7_4__32, linha7_4__31, 
         linha7_4__30, linha7_4__29, linha7_4__28, linha7_4__27, linha7_4__26, 
         linha7_4__25, linha7_4__24, linha7_4__23, linha7_4__22, linha7_4__21, 
         linha7_4__20, linha7_4__19, linha7_4__18, linha7_4__17, linha7_4__16, 
         linha7_4__15, linha7_4__14, linha7_4__13, linha7_4__12, linha7_4__11, 
         linha7_4__10, linha7_4__9, linha7_4__8, linha7_4__7, linha7_4__6, 
         linha7_4__5, linha7_4__4, linha7_4__3, linha7_4__2, linha7_4__1, 
         linha7_4__0, linha7_3__63, linha7_3__62, linha7_3__61, linha7_3__60, 
         linha7_3__59, linha7_3__58, linha7_3__57, linha7_3__56, linha7_3__55, 
         linha7_3__54, linha7_3__53, linha7_3__52, linha7_3__51, linha7_3__50, 
         linha7_3__49, linha7_3__48, linha7_3__47, linha7_3__46, linha7_3__45, 
         linha7_3__44, linha7_3__43, linha7_3__42, linha7_3__41, linha7_3__40, 
         linha7_3__39, linha7_3__38, linha7_3__37, linha7_3__36, linha7_3__35, 
         linha7_3__34, linha7_3__33, linha7_3__32, linha7_3__31, linha7_3__30, 
         linha7_3__29, linha7_3__28, linha7_3__27, linha7_3__26, linha7_3__25, 
         linha7_3__24, linha7_3__23, linha7_3__22, linha7_3__21, linha7_3__20, 
         linha7_3__19, linha7_3__18, linha7_3__17, linha7_3__16, linha7_3__15, 
         linha7_3__14, linha7_3__13, linha7_3__12, linha7_3__11, linha7_3__10, 
         linha7_3__9, linha7_3__8, linha7_3__7, linha7_3__6, linha7_3__5, 
         linha7_3__4, linha7_3__3, linha7_3__2, linha7_3__1, linha7_3__0, 
         linha7_2__63, linha7_2__62, linha7_2__61, linha7_2__60, linha7_2__59, 
         linha7_2__58, linha7_2__57, linha7_2__56, linha7_2__55, linha7_2__54, 
         linha7_2__53, linha7_2__52, linha7_2__51, linha7_2__50, linha7_2__49, 
         linha7_2__48, linha7_2__47, linha7_2__46, linha7_2__45, linha7_2__44, 
         linha7_2__43, linha7_2__42, linha7_2__41, linha7_2__40, linha7_2__39, 
         linha7_2__38, linha7_2__37, linha7_2__36, linha7_2__35, linha7_2__34, 
         linha7_2__33, linha7_2__32, linha7_2__31, linha7_2__30, linha7_2__29, 
         linha7_2__28, linha7_2__27, linha7_2__26, linha7_2__25, linha7_2__24, 
         linha7_2__23, linha7_2__22, linha7_2__21, linha7_2__20, linha7_2__19, 
         linha7_2__18, linha7_2__17, linha7_2__16, linha7_2__15, linha7_2__14, 
         linha7_2__13, linha7_2__12, linha7_2__11, linha7_2__10, linha7_2__9, 
         linha7_2__8, linha7_2__7, linha7_2__6, linha7_2__5, linha7_2__4, 
         linha7_2__3, linha7_2__2, linha7_2__1, linha7_2__0, linha7_1__63, 
         linha7_1__62, linha7_1__61, linha7_1__60, linha7_1__59, linha7_1__58, 
         linha7_1__57, linha7_1__56, linha7_1__55, linha7_1__54, linha7_1__53, 
         linha7_1__52, linha7_1__51, linha7_1__50, linha7_1__49, linha7_1__48, 
         linha7_1__47, linha7_1__46, linha7_1__45, linha7_1__44, linha7_1__43, 
         linha7_1__42, linha7_1__41, linha7_1__40, linha7_1__39, linha7_1__38, 
         linha7_1__37, linha7_1__36, linha7_1__35, linha7_1__34, linha7_1__33, 
         linha7_1__32, linha7_1__31, linha7_1__30, linha7_1__29, linha7_1__28, 
         linha7_1__27, linha7_1__26, linha7_1__25, linha7_1__24, linha7_1__23, 
         linha7_1__22, linha7_1__21, linha7_1__20, linha7_1__19, linha7_1__18, 
         linha7_1__17, linha7_1__16, linha7_1__15, linha7_1__14, linha7_1__13, 
         linha7_1__12, linha7_1__11, linha7_1__10, linha7_1__9, linha7_1__8, 
         linha7_1__7, linha7_1__6, linha7_1__5, linha7_1__4, linha7_1__3, 
         linha7_1__2, linha7_1__1, linha7_1__0, linha6_7__63, linha6_7__62, 
         linha6_7__61, linha6_7__60, linha6_7__59, linha6_7__58, linha6_7__57, 
         linha6_7__56, linha6_7__55, linha6_7__54, linha6_7__53, linha6_7__52, 
         linha6_7__51, linha6_7__50, linha6_7__49, linha6_7__48, linha6_7__47, 
         linha6_7__46, linha6_7__45, linha6_7__44, linha6_7__43, linha6_7__42, 
         linha6_7__41, linha6_7__40, linha6_7__39, linha6_7__38, linha6_7__37, 
         linha6_7__36, linha6_7__35, linha6_7__34, linha6_7__33, linha6_7__32, 
         linha6_7__31, linha6_7__30, linha6_7__29, linha6_7__28, linha6_7__27, 
         linha6_7__26, linha6_7__25, linha6_7__24, linha6_7__23, linha6_7__22, 
         linha6_7__21, linha6_7__20, linha6_7__19, linha6_7__18, linha6_7__17, 
         linha6_7__16, linha6_7__15, linha6_7__14, linha6_7__13, linha6_7__12, 
         linha6_7__11, linha6_7__10, linha6_7__9, linha6_7__8, linha6_7__7, 
         linha6_7__6, linha6_7__5, linha6_7__4, linha6_7__3, linha6_7__2, 
         linha6_7__1, linha6_7__0, linha6_6__63, linha6_6__62, linha6_6__61, 
         linha6_6__60, linha6_6__59, linha6_6__58, linha6_6__57, linha6_6__56, 
         linha6_6__55, linha6_6__54, linha6_6__53, linha6_6__52, linha6_6__51, 
         linha6_6__50, linha6_6__49, linha6_6__48, linha6_6__47, linha6_6__46, 
         linha6_6__45, linha6_6__44, linha6_6__43, linha6_6__42, linha6_6__41, 
         linha6_6__40, linha6_6__39, linha6_6__38, linha6_6__37, linha6_6__36, 
         linha6_6__35, linha6_6__34, linha6_6__33, linha6_6__32, linha6_6__31, 
         linha6_6__30, linha6_6__29, linha6_6__28, linha6_6__27, linha6_6__26, 
         linha6_6__25, linha6_6__24, linha6_6__23, linha6_6__22, linha6_6__21, 
         linha6_6__20, linha6_6__19, linha6_6__18, linha6_6__17, linha6_6__16, 
         linha6_6__15, linha6_6__14, linha6_6__13, linha6_6__12, linha6_6__11, 
         linha6_6__10, linha6_6__9, linha6_6__8, linha6_6__7, linha6_6__6, 
         linha6_6__5, linha6_6__4, linha6_6__3, linha6_6__2, linha6_6__1, 
         linha6_6__0, linha6_5__63, linha6_5__62, linha6_5__61, linha6_5__60, 
         linha6_5__59, linha6_5__58, linha6_5__57, linha6_5__56, linha6_5__55, 
         linha6_5__54, linha6_5__53, linha6_5__52, linha6_5__51, linha6_5__50, 
         linha6_5__49, linha6_5__48, linha6_5__47, linha6_5__46, linha6_5__45, 
         linha6_5__44, linha6_5__43, linha6_5__42, linha6_5__41, linha6_5__40, 
         linha6_5__39, linha6_5__38, linha6_5__37, linha6_5__36, linha6_5__35, 
         linha6_5__34, linha6_5__33, linha6_5__32, linha6_5__31, linha6_5__30, 
         linha6_5__29, linha6_5__28, linha6_5__27, linha6_5__26, linha6_5__25, 
         linha6_5__24, linha6_5__23, linha6_5__22, linha6_5__21, linha6_5__20, 
         linha6_5__19, linha6_5__18, linha6_5__17, linha6_5__16, linha6_5__15, 
         linha6_5__14, linha6_5__13, linha6_5__12, linha6_5__11, linha6_5__10, 
         linha6_5__9, linha6_5__8, linha6_5__7, linha6_5__6, linha6_5__5, 
         linha6_5__4, linha6_5__3, linha6_5__2, linha6_5__1, linha6_5__0, 
         linha6_4__63, linha6_4__62, linha6_4__61, linha6_4__60, linha6_4__59, 
         linha6_4__58, linha6_4__57, linha6_4__56, linha6_4__55, linha6_4__54, 
         linha6_4__53, linha6_4__52, linha6_4__51, linha6_4__50, linha6_4__49, 
         linha6_4__48, linha6_4__47, linha6_4__46, linha6_4__45, linha6_4__44, 
         linha6_4__43, linha6_4__42, linha6_4__41, linha6_4__40, linha6_4__39, 
         linha6_4__38, linha6_4__37, linha6_4__36, linha6_4__35, linha6_4__34, 
         linha6_4__33, linha6_4__32, linha6_4__31, linha6_4__30, linha6_4__29, 
         linha6_4__28, linha6_4__27, linha6_4__26, linha6_4__25, linha6_4__24, 
         linha6_4__23, linha6_4__22, linha6_4__21, linha6_4__20, linha6_4__19, 
         linha6_4__18, linha6_4__17, linha6_4__16, linha6_4__15, linha6_4__14, 
         linha6_4__13, linha6_4__12, linha6_4__11, linha6_4__10, linha6_4__9, 
         linha6_4__8, linha6_4__7, linha6_4__6, linha6_4__5, linha6_4__4, 
         linha6_4__3, linha6_4__2, linha6_4__1, linha6_4__0, linha6_3__63, 
         linha6_3__62, linha6_3__61, linha6_3__60, linha6_3__59, linha6_3__58, 
         linha6_3__57, linha6_3__56, linha6_3__55, linha6_3__54, linha6_3__53, 
         linha6_3__52, linha6_3__51, linha6_3__50, linha6_3__49, linha6_3__48, 
         linha6_3__47, linha6_3__46, linha6_3__45, linha6_3__44, linha6_3__43, 
         linha6_3__42, linha6_3__41, linha6_3__40, linha6_3__39, linha6_3__38, 
         linha6_3__37, linha6_3__36, linha6_3__35, linha6_3__34, linha6_3__33, 
         linha6_3__32, linha6_3__31, linha6_3__30, linha6_3__29, linha6_3__28, 
         linha6_3__27, linha6_3__26, linha6_3__25, linha6_3__24, linha6_3__23, 
         linha6_3__22, linha6_3__21, linha6_3__20, linha6_3__19, linha6_3__18, 
         linha6_3__17, linha6_3__16, linha6_3__15, linha6_3__14, linha6_3__13, 
         linha6_3__12, linha6_3__11, linha6_3__10, linha6_3__9, linha6_3__8, 
         linha6_3__7, linha6_3__6, linha6_3__5, linha6_3__4, linha6_3__3, 
         linha6_3__2, linha6_3__1, linha6_3__0, linha6_2__63, linha6_2__62, 
         linha6_2__61, linha6_2__60, linha6_2__59, linha6_2__58, linha6_2__57, 
         linha6_2__56, linha6_2__55, linha6_2__54, linha6_2__53, linha6_2__52, 
         linha6_2__51, linha6_2__50, linha6_2__49, linha6_2__48, linha6_2__47, 
         linha6_2__46, linha6_2__45, linha6_2__44, linha6_2__43, linha6_2__42, 
         linha6_2__41, linha6_2__40, linha6_2__39, linha6_2__38, linha6_2__37, 
         linha6_2__36, linha6_2__35, linha6_2__34, linha6_2__33, linha6_2__32, 
         linha6_2__31, linha6_2__30, linha6_2__29, linha6_2__28, linha6_2__27, 
         linha6_2__26, linha6_2__25, linha6_2__24, linha6_2__23, linha6_2__22, 
         linha6_2__21, linha6_2__20, linha6_2__19, linha6_2__18, linha6_2__17, 
         linha6_2__16, linha6_2__15, linha6_2__14, linha6_2__13, linha6_2__12, 
         linha6_2__11, linha6_2__10, linha6_2__9, linha6_2__8, linha6_2__7, 
         linha6_2__6, linha6_2__5, linha6_2__4, linha6_2__3, linha6_2__2, 
         linha6_2__1, linha6_2__0, linha6_1__63, linha6_1__62, linha6_1__61, 
         linha6_1__60, linha6_1__59, linha6_1__58, linha6_1__57, linha6_1__56, 
         linha6_1__55, linha6_1__54, linha6_1__53, linha6_1__52, linha6_1__51, 
         linha6_1__50, linha6_1__49, linha6_1__48, linha6_1__47, linha6_1__46, 
         linha6_1__45, linha6_1__44, linha6_1__43, linha6_1__42, linha6_1__41, 
         linha6_1__40, linha6_1__39, linha6_1__38, linha6_1__37, linha6_1__36, 
         linha6_1__35, linha6_1__34, linha6_1__33, linha6_1__32, linha6_1__31, 
         linha6_1__30, linha6_1__29, linha6_1__28, linha6_1__27, linha6_1__26, 
         linha6_1__25, linha6_1__24, linha6_1__23, linha6_1__22, linha6_1__21, 
         linha6_1__20, linha6_1__19, linha6_1__18, linha6_1__17, linha6_1__16, 
         linha6_1__15, linha6_1__14, linha6_1__13, linha6_1__12, linha6_1__11, 
         linha6_1__10, linha6_1__9, linha6_1__8, linha6_1__7, linha6_1__6, 
         linha6_1__5, linha6_1__4, linha6_1__3, linha6_1__2, linha6_1__1, 
         linha6_1__0, linha5_7__63, linha5_7__62, linha5_7__61, linha5_7__60, 
         linha5_7__59, linha5_7__58, linha5_7__57, linha5_7__56, linha5_7__55, 
         linha5_7__54, linha5_7__53, linha5_7__52, linha5_7__51, linha5_7__50, 
         linha5_7__49, linha5_7__48, linha5_7__47, linha5_7__46, linha5_7__45, 
         linha5_7__44, linha5_7__43, linha5_7__42, linha5_7__41, linha5_7__40, 
         linha5_7__39, linha5_7__38, linha5_7__37, linha5_7__36, linha5_7__35, 
         linha5_7__34, linha5_7__33, linha5_7__32, linha5_7__31, linha5_7__30, 
         linha5_7__29, linha5_7__28, linha5_7__27, linha5_7__26, linha5_7__25, 
         linha5_7__24, linha5_7__23, linha5_7__22, linha5_7__21, linha5_7__20, 
         linha5_7__19, linha5_7__18, linha5_7__17, linha5_7__16, linha5_7__15, 
         linha5_7__14, linha5_7__13, linha5_7__12, linha5_7__11, linha5_7__10, 
         linha5_7__9, linha5_7__8, linha5_7__7, linha5_7__6, linha5_7__5, 
         linha5_7__4, linha5_7__3, linha5_7__2, linha5_7__1, linha5_7__0, 
         linha5_6__63, linha5_6__62, linha5_6__61, linha5_6__60, linha5_6__59, 
         linha5_6__58, linha5_6__57, linha5_6__56, linha5_6__55, linha5_6__54, 
         linha5_6__53, linha5_6__52, linha5_6__51, linha5_6__50, linha5_6__49, 
         linha5_6__48, linha5_6__47, linha5_6__46, linha5_6__45, linha5_6__44, 
         linha5_6__43, linha5_6__42, linha5_6__41, linha5_6__40, linha5_6__39, 
         linha5_6__38, linha5_6__37, linha5_6__36, linha5_6__35, linha5_6__34, 
         linha5_6__33, linha5_6__32, linha5_6__31, linha5_6__30, linha5_6__29, 
         linha5_6__28, linha5_6__27, linha5_6__26, linha5_6__25, linha5_6__24, 
         linha5_6__23, linha5_6__22, linha5_6__21, linha5_6__20, linha5_6__19, 
         linha5_6__18, linha5_6__17, linha5_6__16, linha5_6__15, linha5_6__14, 
         linha5_6__13, linha5_6__12, linha5_6__11, linha5_6__10, linha5_6__9, 
         linha5_6__8, linha5_6__7, linha5_6__6, linha5_6__5, linha5_6__4, 
         linha5_6__3, linha5_6__2, linha5_6__1, linha5_6__0, linha5_5__63, 
         linha5_5__62, linha5_5__61, linha5_5__60, linha5_5__59, linha5_5__58, 
         linha5_5__57, linha5_5__56, linha5_5__55, linha5_5__54, linha5_5__53, 
         linha5_5__52, linha5_5__51, linha5_5__50, linha5_5__49, linha5_5__48, 
         linha5_5__47, linha5_5__46, linha5_5__45, linha5_5__44, linha5_5__43, 
         linha5_5__42, linha5_5__41, linha5_5__40, linha5_5__39, linha5_5__38, 
         linha5_5__37, linha5_5__36, linha5_5__35, linha5_5__34, linha5_5__33, 
         linha5_5__32, linha5_5__31, linha5_5__30, linha5_5__29, linha5_5__28, 
         linha5_5__27, linha5_5__26, linha5_5__25, linha5_5__24, linha5_5__23, 
         linha5_5__22, linha5_5__21, linha5_5__20, linha5_5__19, linha5_5__18, 
         linha5_5__17, linha5_5__16, linha5_5__15, linha5_5__14, linha5_5__13, 
         linha5_5__12, linha5_5__11, linha5_5__10, linha5_5__9, linha5_5__8, 
         linha5_5__7, linha5_5__6, linha5_5__5, linha5_5__4, linha5_5__3, 
         linha5_5__2, linha5_5__1, linha5_5__0, linha5_4__63, linha5_4__62, 
         linha5_4__61, linha5_4__60, linha5_4__59, linha5_4__58, linha5_4__57, 
         linha5_4__56, linha5_4__55, linha5_4__54, linha5_4__53, linha5_4__52, 
         linha5_4__51, linha5_4__50, linha5_4__49, linha5_4__48, linha5_4__47, 
         linha5_4__46, linha5_4__45, linha5_4__44, linha5_4__43, linha5_4__42, 
         linha5_4__41, linha5_4__40, linha5_4__39, linha5_4__38, linha5_4__37, 
         linha5_4__36, linha5_4__35, linha5_4__34, linha5_4__33, linha5_4__32, 
         linha5_4__31, linha5_4__30, linha5_4__29, linha5_4__28, linha5_4__27, 
         linha5_4__26, linha5_4__25, linha5_4__24, linha5_4__23, linha5_4__22, 
         linha5_4__21, linha5_4__20, linha5_4__19, linha5_4__18, linha5_4__17, 
         linha5_4__16, linha5_4__15, linha5_4__14, linha5_4__13, linha5_4__12, 
         linha5_4__11, linha5_4__10, linha5_4__9, linha5_4__8, linha5_4__7, 
         linha5_4__6, linha5_4__5, linha5_4__4, linha5_4__3, linha5_4__2, 
         linha5_4__1, linha5_4__0, linha5_3__63, linha5_3__62, linha5_3__61, 
         linha5_3__60, linha5_3__59, linha5_3__58, linha5_3__57, linha5_3__56, 
         linha5_3__55, linha5_3__54, linha5_3__53, linha5_3__52, linha5_3__51, 
         linha5_3__50, linha5_3__49, linha5_3__48, linha5_3__47, linha5_3__46, 
         linha5_3__45, linha5_3__44, linha5_3__43, linha5_3__42, linha5_3__41, 
         linha5_3__40, linha5_3__39, linha5_3__38, linha5_3__37, linha5_3__36, 
         linha5_3__35, linha5_3__34, linha5_3__33, linha5_3__32, linha5_3__31, 
         linha5_3__30, linha5_3__29, linha5_3__28, linha5_3__27, linha5_3__26, 
         linha5_3__25, linha5_3__24, linha5_3__23, linha5_3__22, linha5_3__21, 
         linha5_3__20, linha5_3__19, linha5_3__18, linha5_3__17, linha5_3__16, 
         linha5_3__15, linha5_3__14, linha5_3__13, linha5_3__12, linha5_3__11, 
         linha5_3__10, linha5_3__9, linha5_3__8, linha5_3__7, linha5_3__6, 
         linha5_3__5, linha5_3__4, linha5_3__3, linha5_3__2, linha5_3__1, 
         linha5_3__0, linha5_2__63, linha5_2__62, linha5_2__61, linha5_2__60, 
         linha5_2__59, linha5_2__58, linha5_2__57, linha5_2__56, linha5_2__55, 
         linha5_2__54, linha5_2__53, linha5_2__52, linha5_2__51, linha5_2__50, 
         linha5_2__49, linha5_2__48, linha5_2__47, linha5_2__46, linha5_2__45, 
         linha5_2__44, linha5_2__43, linha5_2__42, linha5_2__41, linha5_2__40, 
         linha5_2__39, linha5_2__38, linha5_2__37, linha5_2__36, linha5_2__35, 
         linha5_2__34, linha5_2__33, linha5_2__32, linha5_2__31, linha5_2__30, 
         linha5_2__29, linha5_2__28, linha5_2__27, linha5_2__26, linha5_2__25, 
         linha5_2__24, linha5_2__23, linha5_2__22, linha5_2__21, linha5_2__20, 
         linha5_2__19, linha5_2__18, linha5_2__17, linha5_2__16, linha5_2__15, 
         linha5_2__14, linha5_2__13, linha5_2__12, linha5_2__11, linha5_2__10, 
         linha5_2__9, linha5_2__8, linha5_2__7, linha5_2__6, linha5_2__5, 
         linha5_2__4, linha5_2__3, linha5_2__2, linha5_2__1, linha5_2__0, 
         linha5_1__63, linha5_1__62, linha5_1__61, linha5_1__60, linha5_1__59, 
         linha5_1__58, linha5_1__57, linha5_1__56, linha5_1__55, linha5_1__54, 
         linha5_1__53, linha5_1__52, linha5_1__51, linha5_1__50, linha5_1__49, 
         linha5_1__48, linha5_1__47, linha5_1__46, linha5_1__45, linha5_1__44, 
         linha5_1__43, linha5_1__42, linha5_1__41, linha5_1__40, linha5_1__39, 
         linha5_1__38, linha5_1__37, linha5_1__36, linha5_1__35, linha5_1__34, 
         linha5_1__33, linha5_1__32, linha5_1__31, linha5_1__30, linha5_1__29, 
         linha5_1__28, linha5_1__27, linha5_1__26, linha5_1__25, linha5_1__24, 
         linha5_1__23, linha5_1__22, linha5_1__21, linha5_1__20, linha5_1__19, 
         linha5_1__18, linha5_1__17, linha5_1__16, linha5_1__15, linha5_1__14, 
         linha5_1__13, linha5_1__12, linha5_1__11, linha5_1__10, linha5_1__9, 
         linha5_1__8, linha5_1__7, linha5_1__6, linha5_1__5, linha5_1__4, 
         linha5_1__3, linha5_1__2, linha5_1__1, linha5_1__0, linha4_7__63, 
         linha4_7__62, linha4_7__61, linha4_7__60, linha4_7__59, linha4_7__58, 
         linha4_7__57, linha4_7__56, linha4_7__55, linha4_7__54, linha4_7__53, 
         linha4_7__52, linha4_7__51, linha4_7__50, linha4_7__49, linha4_7__48, 
         linha4_7__47, linha4_7__46, linha4_7__45, linha4_7__44, linha4_7__43, 
         linha4_7__42, linha4_7__41, linha4_7__40, linha4_7__39, linha4_7__38, 
         linha4_7__37, linha4_7__36, linha4_7__35, linha4_7__34, linha4_7__33, 
         linha4_7__32, linha4_7__31, linha4_7__30, linha4_7__29, linha4_7__28, 
         linha4_7__27, linha4_7__26, linha4_7__25, linha4_7__24, linha4_7__23, 
         linha4_7__22, linha4_7__21, linha4_7__20, linha4_7__19, linha4_7__18, 
         linha4_7__17, linha4_7__16, linha4_7__15, linha4_7__14, linha4_7__13, 
         linha4_7__12, linha4_7__11, linha4_7__10, linha4_7__9, linha4_7__8, 
         linha4_7__7, linha4_7__6, linha4_7__5, linha4_7__4, linha4_7__3, 
         linha4_7__2, linha4_7__1, linha4_7__0, linha4_6__63, linha4_6__62, 
         linha4_6__61, linha4_6__60, linha4_6__59, linha4_6__58, linha4_6__57, 
         linha4_6__56, linha4_6__55, linha4_6__54, linha4_6__53, linha4_6__52, 
         linha4_6__51, linha4_6__50, linha4_6__49, linha4_6__48, linha4_6__47, 
         linha4_6__46, linha4_6__45, linha4_6__44, linha4_6__43, linha4_6__42, 
         linha4_6__41, linha4_6__40, linha4_6__39, linha4_6__38, linha4_6__37, 
         linha4_6__36, linha4_6__35, linha4_6__34, linha4_6__33, linha4_6__32, 
         linha4_6__31, linha4_6__30, linha4_6__29, linha4_6__28, linha4_6__27, 
         linha4_6__26, linha4_6__25, linha4_6__24, linha4_6__23, linha4_6__22, 
         linha4_6__21, linha4_6__20, linha4_6__19, linha4_6__18, linha4_6__17, 
         linha4_6__16, linha4_6__15, linha4_6__14, linha4_6__13, linha4_6__12, 
         linha4_6__11, linha4_6__10, linha4_6__9, linha4_6__8, linha4_6__7, 
         linha4_6__6, linha4_6__5, linha4_6__4, linha4_6__3, linha4_6__2, 
         linha4_6__1, linha4_6__0, linha4_5__63, linha4_5__62, linha4_5__61, 
         linha4_5__60, linha4_5__59, linha4_5__58, linha4_5__57, linha4_5__56, 
         linha4_5__55, linha4_5__54, linha4_5__53, linha4_5__52, linha4_5__51, 
         linha4_5__50, linha4_5__49, linha4_5__48, linha4_5__47, linha4_5__46, 
         linha4_5__45, linha4_5__44, linha4_5__43, linha4_5__42, linha4_5__41, 
         linha4_5__40, linha4_5__39, linha4_5__38, linha4_5__37, linha4_5__36, 
         linha4_5__35, linha4_5__34, linha4_5__33, linha4_5__32, linha4_5__31, 
         linha4_5__30, linha4_5__29, linha4_5__28, linha4_5__27, linha4_5__26, 
         linha4_5__25, linha4_5__24, linha4_5__23, linha4_5__22, linha4_5__21, 
         linha4_5__20, linha4_5__19, linha4_5__18, linha4_5__17, linha4_5__16, 
         linha4_5__15, linha4_5__14, linha4_5__13, linha4_5__12, linha4_5__11, 
         linha4_5__10, linha4_5__9, linha4_5__8, linha4_5__7, linha4_5__6, 
         linha4_5__5, linha4_5__4, linha4_5__3, linha4_5__2, linha4_5__1, 
         linha4_5__0, linha4_4__63, linha4_4__62, linha4_4__61, linha4_4__60, 
         linha4_4__59, linha4_4__58, linha4_4__57, linha4_4__56, linha4_4__55, 
         linha4_4__54, linha4_4__53, linha4_4__52, linha4_4__51, linha4_4__50, 
         linha4_4__49, linha4_4__48, linha4_4__47, linha4_4__46, linha4_4__45, 
         linha4_4__44, linha4_4__43, linha4_4__42, linha4_4__41, linha4_4__40, 
         linha4_4__39, linha4_4__38, linha4_4__37, linha4_4__36, linha4_4__35, 
         linha4_4__34, linha4_4__33, linha4_4__32, linha4_4__31, linha4_4__30, 
         linha4_4__29, linha4_4__28, linha4_4__27, linha4_4__26, linha4_4__25, 
         linha4_4__24, linha4_4__23, linha4_4__22, linha4_4__21, linha4_4__20, 
         linha4_4__19, linha4_4__18, linha4_4__17, linha4_4__16, linha4_4__15, 
         linha4_4__14, linha4_4__13, linha4_4__12, linha4_4__11, linha4_4__10, 
         linha4_4__9, linha4_4__8, linha4_4__7, linha4_4__6, linha4_4__5, 
         linha4_4__4, linha4_4__3, linha4_4__2, linha4_4__1, linha4_4__0, 
         linha4_3__63, linha4_3__62, linha4_3__61, linha4_3__60, linha4_3__59, 
         linha4_3__58, linha4_3__57, linha4_3__56, linha4_3__55, linha4_3__54, 
         linha4_3__53, linha4_3__52, linha4_3__51, linha4_3__50, linha4_3__49, 
         linha4_3__48, linha4_3__47, linha4_3__46, linha4_3__45, linha4_3__44, 
         linha4_3__43, linha4_3__42, linha4_3__41, linha4_3__40, linha4_3__39, 
         linha4_3__38, linha4_3__37, linha4_3__36, linha4_3__35, linha4_3__34, 
         linha4_3__33, linha4_3__32, linha4_3__31, linha4_3__30, linha4_3__29, 
         linha4_3__28, linha4_3__27, linha4_3__26, linha4_3__25, linha4_3__24, 
         linha4_3__23, linha4_3__22, linha4_3__21, linha4_3__20, linha4_3__19, 
         linha4_3__18, linha4_3__17, linha4_3__16, linha4_3__15, linha4_3__14, 
         linha4_3__13, linha4_3__12, linha4_3__11, linha4_3__10, linha4_3__9, 
         linha4_3__8, linha4_3__7, linha4_3__6, linha4_3__5, linha4_3__4, 
         linha4_3__3, linha4_3__2, linha4_3__1, linha4_3__0, linha4_2__63, 
         linha4_2__62, linha4_2__61, linha4_2__60, linha4_2__59, linha4_2__58, 
         linha4_2__57, linha4_2__56, linha4_2__55, linha4_2__54, linha4_2__53, 
         linha4_2__52, linha4_2__51, linha4_2__50, linha4_2__49, linha4_2__48, 
         linha4_2__47, linha4_2__46, linha4_2__45, linha4_2__44, linha4_2__43, 
         linha4_2__42, linha4_2__41, linha4_2__40, linha4_2__39, linha4_2__38, 
         linha4_2__37, linha4_2__36, linha4_2__35, linha4_2__34, linha4_2__33, 
         linha4_2__32, linha4_2__31, linha4_2__30, linha4_2__29, linha4_2__28, 
         linha4_2__27, linha4_2__26, linha4_2__25, linha4_2__24, linha4_2__23, 
         linha4_2__22, linha4_2__21, linha4_2__20, linha4_2__19, linha4_2__18, 
         linha4_2__17, linha4_2__16, linha4_2__15, linha4_2__14, linha4_2__13, 
         linha4_2__12, linha4_2__11, linha4_2__10, linha4_2__9, linha4_2__8, 
         linha4_2__7, linha4_2__6, linha4_2__5, linha4_2__4, linha4_2__3, 
         linha4_2__2, linha4_2__1, linha4_2__0, linha4_1__63, linha4_1__62, 
         linha4_1__61, linha4_1__60, linha4_1__59, linha4_1__58, linha4_1__57, 
         linha4_1__56, linha4_1__55, linha4_1__54, linha4_1__53, linha4_1__52, 
         linha4_1__51, linha4_1__50, linha4_1__49, linha4_1__48, linha4_1__47, 
         linha4_1__46, linha4_1__45, linha4_1__44, linha4_1__43, linha4_1__42, 
         linha4_1__41, linha4_1__40, linha4_1__39, linha4_1__38, linha4_1__37, 
         linha4_1__36, linha4_1__35, linha4_1__34, linha4_1__33, linha4_1__32, 
         linha4_1__31, linha4_1__30, linha4_1__29, linha4_1__28, linha4_1__27, 
         linha4_1__26, linha4_1__25, linha4_1__24, linha4_1__23, linha4_1__22, 
         linha4_1__21, linha4_1__20, linha4_1__19, linha4_1__18, linha4_1__17, 
         linha4_1__16, linha4_1__15, linha4_1__14, linha4_1__13, linha4_1__12, 
         linha4_1__11, linha4_1__10, linha4_1__9, linha4_1__8, linha4_1__7, 
         linha4_1__6, linha4_1__5, linha4_1__4, linha4_1__3, linha4_1__2, 
         linha4_1__1, linha4_1__0, linha3_7__63, linha3_7__62, linha3_7__61, 
         linha3_7__60, linha3_7__59, linha3_7__58, linha3_7__57, linha3_7__56, 
         linha3_7__55, linha3_7__54, linha3_7__53, linha3_7__52, linha3_7__51, 
         linha3_7__50, linha3_7__49, linha3_7__48, linha3_7__47, linha3_7__46, 
         linha3_7__45, linha3_7__44, linha3_7__43, linha3_7__42, linha3_7__41, 
         linha3_7__40, linha3_7__39, linha3_7__38, linha3_7__37, linha3_7__36, 
         linha3_7__35, linha3_7__34, linha3_7__33, linha3_7__32, linha3_7__31, 
         linha3_7__30, linha3_7__29, linha3_7__28, linha3_7__27, linha3_7__26, 
         linha3_7__25, linha3_7__24, linha3_7__23, linha3_7__22, linha3_7__21, 
         linha3_7__20, linha3_7__19, linha3_7__18, linha3_7__17, linha3_7__16, 
         linha3_7__15, linha3_7__14, linha3_7__13, linha3_7__12, linha3_7__11, 
         linha3_7__10, linha3_7__9, linha3_7__8, linha3_7__7, linha3_7__6, 
         linha3_7__5, linha3_7__4, linha3_7__3, linha3_7__2, linha3_7__1, 
         linha3_7__0, linha3_6__63, linha3_6__62, linha3_6__61, linha3_6__60, 
         linha3_6__59, linha3_6__58, linha3_6__57, linha3_6__56, linha3_6__55, 
         linha3_6__54, linha3_6__53, linha3_6__52, linha3_6__51, linha3_6__50, 
         linha3_6__49, linha3_6__48, linha3_6__47, linha3_6__46, linha3_6__45, 
         linha3_6__44, linha3_6__43, linha3_6__42, linha3_6__41, linha3_6__40, 
         linha3_6__39, linha3_6__38, linha3_6__37, linha3_6__36, linha3_6__35, 
         linha3_6__34, linha3_6__33, linha3_6__32, linha3_6__31, linha3_6__30, 
         linha3_6__29, linha3_6__28, linha3_6__27, linha3_6__26, linha3_6__25, 
         linha3_6__24, linha3_6__23, linha3_6__22, linha3_6__21, linha3_6__20, 
         linha3_6__19, linha3_6__18, linha3_6__17, linha3_6__16, linha3_6__15, 
         linha3_6__14, linha3_6__13, linha3_6__12, linha3_6__11, linha3_6__10, 
         linha3_6__9, linha3_6__8, linha3_6__7, linha3_6__6, linha3_6__5, 
         linha3_6__4, linha3_6__3, linha3_6__2, linha3_6__1, linha3_6__0, 
         linha3_5__63, linha3_5__62, linha3_5__61, linha3_5__60, linha3_5__59, 
         linha3_5__58, linha3_5__57, linha3_5__56, linha3_5__55, linha3_5__54, 
         linha3_5__53, linha3_5__52, linha3_5__51, linha3_5__50, linha3_5__49, 
         linha3_5__48, linha3_5__47, linha3_5__46, linha3_5__45, linha3_5__44, 
         linha3_5__43, linha3_5__42, linha3_5__41, linha3_5__40, linha3_5__39, 
         linha3_5__38, linha3_5__37, linha3_5__36, linha3_5__35, linha3_5__34, 
         linha3_5__33, linha3_5__32, linha3_5__31, linha3_5__30, linha3_5__29, 
         linha3_5__28, linha3_5__27, linha3_5__26, linha3_5__25, linha3_5__24, 
         linha3_5__23, linha3_5__22, linha3_5__21, linha3_5__20, linha3_5__19, 
         linha3_5__18, linha3_5__17, linha3_5__16, linha3_5__15, linha3_5__14, 
         linha3_5__13, linha3_5__12, linha3_5__11, linha3_5__10, linha3_5__9, 
         linha3_5__8, linha3_5__7, linha3_5__6, linha3_5__5, linha3_5__4, 
         linha3_5__3, linha3_5__2, linha3_5__1, linha3_5__0, linha3_4__63, 
         linha3_4__62, linha3_4__61, linha3_4__60, linha3_4__59, linha3_4__58, 
         linha3_4__57, linha3_4__56, linha3_4__55, linha3_4__54, linha3_4__53, 
         linha3_4__52, linha3_4__51, linha3_4__50, linha3_4__49, linha3_4__48, 
         linha3_4__47, linha3_4__46, linha3_4__45, linha3_4__44, linha3_4__43, 
         linha3_4__42, linha3_4__41, linha3_4__40, linha3_4__39, linha3_4__38, 
         linha3_4__37, linha3_4__36, linha3_4__35, linha3_4__34, linha3_4__33, 
         linha3_4__32, linha3_4__31, linha3_4__30, linha3_4__29, linha3_4__28, 
         linha3_4__27, linha3_4__26, linha3_4__25, linha3_4__24, linha3_4__23, 
         linha3_4__22, linha3_4__21, linha3_4__20, linha3_4__19, linha3_4__18, 
         linha3_4__17, linha3_4__16, linha3_4__15, linha3_4__14, linha3_4__13, 
         linha3_4__12, linha3_4__11, linha3_4__10, linha3_4__9, linha3_4__8, 
         linha3_4__7, linha3_4__6, linha3_4__5, linha3_4__4, linha3_4__3, 
         linha3_4__2, linha3_4__1, linha3_4__0, linha3_3__63, linha3_3__62, 
         linha3_3__61, linha3_3__60, linha3_3__59, linha3_3__58, linha3_3__57, 
         linha3_3__56, linha3_3__55, linha3_3__54, linha3_3__53, linha3_3__52, 
         linha3_3__51, linha3_3__50, linha3_3__49, linha3_3__48, linha3_3__47, 
         linha3_3__46, linha3_3__45, linha3_3__44, linha3_3__43, linha3_3__42, 
         linha3_3__41, linha3_3__40, linha3_3__39, linha3_3__38, linha3_3__37, 
         linha3_3__36, linha3_3__35, linha3_3__34, linha3_3__33, linha3_3__32, 
         linha3_3__31, linha3_3__30, linha3_3__29, linha3_3__28, linha3_3__27, 
         linha3_3__26, linha3_3__25, linha3_3__24, linha3_3__23, linha3_3__22, 
         linha3_3__21, linha3_3__20, linha3_3__19, linha3_3__18, linha3_3__17, 
         linha3_3__16, linha3_3__15, linha3_3__14, linha3_3__13, linha3_3__12, 
         linha3_3__11, linha3_3__10, linha3_3__9, linha3_3__8, linha3_3__7, 
         linha3_3__6, linha3_3__5, linha3_3__4, linha3_3__3, linha3_3__2, 
         linha3_3__1, linha3_3__0, linha3_2__63, linha3_2__62, linha3_2__61, 
         linha3_2__60, linha3_2__59, linha3_2__58, linha3_2__57, linha3_2__56, 
         linha3_2__55, linha3_2__54, linha3_2__53, linha3_2__52, linha3_2__51, 
         linha3_2__50, linha3_2__49, linha3_2__48, linha3_2__47, linha3_2__46, 
         linha3_2__45, linha3_2__44, linha3_2__43, linha3_2__42, linha3_2__41, 
         linha3_2__40, linha3_2__39, linha3_2__38, linha3_2__37, linha3_2__36, 
         linha3_2__35, linha3_2__34, linha3_2__33, linha3_2__32, linha3_2__31, 
         linha3_2__30, linha3_2__29, linha3_2__28, linha3_2__27, linha3_2__26, 
         linha3_2__25, linha3_2__24, linha3_2__23, linha3_2__22, linha3_2__21, 
         linha3_2__20, linha3_2__19, linha3_2__18, linha3_2__17, linha3_2__16, 
         linha3_2__15, linha3_2__14, linha3_2__13, linha3_2__12, linha3_2__11, 
         linha3_2__10, linha3_2__9, linha3_2__8, linha3_2__7, linha3_2__6, 
         linha3_2__5, linha3_2__4, linha3_2__3, linha3_2__2, linha3_2__1, 
         linha3_2__0, linha3_1__63, linha3_1__62, linha3_1__61, linha3_1__60, 
         linha3_1__59, linha3_1__58, linha3_1__57, linha3_1__56, linha3_1__55, 
         linha3_1__54, linha3_1__53, linha3_1__52, linha3_1__51, linha3_1__50, 
         linha3_1__49, linha3_1__48, linha3_1__47, linha3_1__46, linha3_1__45, 
         linha3_1__44, linha3_1__43, linha3_1__42, linha3_1__41, linha3_1__40, 
         linha3_1__39, linha3_1__38, linha3_1__37, linha3_1__36, linha3_1__35, 
         linha3_1__34, linha3_1__33, linha3_1__32, linha3_1__31, linha3_1__30, 
         linha3_1__29, linha3_1__28, linha3_1__27, linha3_1__26, linha3_1__25, 
         linha3_1__24, linha3_1__23, linha3_1__22, linha3_1__21, linha3_1__20, 
         linha3_1__19, linha3_1__18, linha3_1__17, linha3_1__16, linha3_1__15, 
         linha3_1__14, linha3_1__13, linha3_1__12, linha3_1__11, linha3_1__10, 
         linha3_1__9, linha3_1__8, linha3_1__7, linha3_1__6, linha3_1__5, 
         linha3_1__4, linha3_1__3, linha3_1__2, linha3_1__1, linha3_1__0, 
         linha2_7__63, linha2_7__62, linha2_7__61, linha2_7__60, linha2_7__59, 
         linha2_7__58, linha2_7__57, linha2_7__56, linha2_7__55, linha2_7__54, 
         linha2_7__53, linha2_7__52, linha2_7__51, linha2_7__50, linha2_7__49, 
         linha2_7__48, linha2_7__47, linha2_7__46, linha2_7__45, linha2_7__44, 
         linha2_7__43, linha2_7__42, linha2_7__41, linha2_7__40, linha2_7__39, 
         linha2_7__38, linha2_7__37, linha2_7__36, linha2_7__35, linha2_7__34, 
         linha2_7__33, linha2_7__32, linha2_7__31, linha2_7__30, linha2_7__29, 
         linha2_7__28, linha2_7__27, linha2_7__26, linha2_7__25, linha2_7__24, 
         linha2_7__23, linha2_7__22, linha2_7__21, linha2_7__20, linha2_7__19, 
         linha2_7__18, linha2_7__17, linha2_7__16, linha2_7__15, linha2_7__14, 
         linha2_7__13, linha2_7__12, linha2_7__11, linha2_7__10, linha2_7__9, 
         linha2_7__8, linha2_7__7, linha2_7__6, linha2_7__5, linha2_7__4, 
         linha2_7__3, linha2_7__2, linha2_7__1, linha2_7__0, linha2_6__63, 
         linha2_6__62, linha2_6__61, linha2_6__60, linha2_6__59, linha2_6__58, 
         linha2_6__57, linha2_6__56, linha2_6__55, linha2_6__54, linha2_6__53, 
         linha2_6__52, linha2_6__51, linha2_6__50, linha2_6__49, linha2_6__48, 
         linha2_6__47, linha2_6__46, linha2_6__45, linha2_6__44, linha2_6__43, 
         linha2_6__42, linha2_6__41, linha2_6__40, linha2_6__39, linha2_6__38, 
         linha2_6__37, linha2_6__36, linha2_6__35, linha2_6__34, linha2_6__33, 
         linha2_6__32, linha2_6__31, linha2_6__30, linha2_6__29, linha2_6__28, 
         linha2_6__27, linha2_6__26, linha2_6__25, linha2_6__24, linha2_6__23, 
         linha2_6__22, linha2_6__21, linha2_6__20, linha2_6__19, linha2_6__18, 
         linha2_6__17, linha2_6__16, linha2_6__15, linha2_6__14, linha2_6__13, 
         linha2_6__12, linha2_6__11, linha2_6__10, linha2_6__9, linha2_6__8, 
         linha2_6__7, linha2_6__6, linha2_6__5, linha2_6__4, linha2_6__3, 
         linha2_6__2, linha2_6__1, linha2_6__0, linha2_5__63, linha2_5__62, 
         linha2_5__61, linha2_5__60, linha2_5__59, linha2_5__58, linha2_5__57, 
         linha2_5__56, linha2_5__55, linha2_5__54, linha2_5__53, linha2_5__52, 
         linha2_5__51, linha2_5__50, linha2_5__49, linha2_5__48, linha2_5__47, 
         linha2_5__46, linha2_5__45, linha2_5__44, linha2_5__43, linha2_5__42, 
         linha2_5__41, linha2_5__40, linha2_5__39, linha2_5__38, linha2_5__37, 
         linha2_5__36, linha2_5__35, linha2_5__34, linha2_5__33, linha2_5__32, 
         linha2_5__31, linha2_5__30, linha2_5__29, linha2_5__28, linha2_5__27, 
         linha2_5__26, linha2_5__25, linha2_5__24, linha2_5__23, linha2_5__22, 
         linha2_5__21, linha2_5__20, linha2_5__19, linha2_5__18, linha2_5__17, 
         linha2_5__16, linha2_5__15, linha2_5__14, linha2_5__13, linha2_5__12, 
         linha2_5__11, linha2_5__10, linha2_5__9, linha2_5__8, linha2_5__7, 
         linha2_5__6, linha2_5__5, linha2_5__4, linha2_5__3, linha2_5__2, 
         linha2_5__1, linha2_5__0, linha2_4__63, linha2_4__62, linha2_4__61, 
         linha2_4__60, linha2_4__59, linha2_4__58, linha2_4__57, linha2_4__56, 
         linha2_4__55, linha2_4__54, linha2_4__53, linha2_4__52, linha2_4__51, 
         linha2_4__50, linha2_4__49, linha2_4__48, linha2_4__47, linha2_4__46, 
         linha2_4__45, linha2_4__44, linha2_4__43, linha2_4__42, linha2_4__41, 
         linha2_4__40, linha2_4__39, linha2_4__38, linha2_4__37, linha2_4__36, 
         linha2_4__35, linha2_4__34, linha2_4__33, linha2_4__32, linha2_4__31, 
         linha2_4__30, linha2_4__29, linha2_4__28, linha2_4__27, linha2_4__26, 
         linha2_4__25, linha2_4__24, linha2_4__23, linha2_4__22, linha2_4__21, 
         linha2_4__20, linha2_4__19, linha2_4__18, linha2_4__17, linha2_4__16, 
         linha2_4__15, linha2_4__14, linha2_4__13, linha2_4__12, linha2_4__11, 
         linha2_4__10, linha2_4__9, linha2_4__8, linha2_4__7, linha2_4__6, 
         linha2_4__5, linha2_4__4, linha2_4__3, linha2_4__2, linha2_4__1, 
         linha2_4__0, linha2_3__63, linha2_3__62, linha2_3__61, linha2_3__60, 
         linha2_3__59, linha2_3__58, linha2_3__57, linha2_3__56, linha2_3__55, 
         linha2_3__54, linha2_3__53, linha2_3__52, linha2_3__51, linha2_3__50, 
         linha2_3__49, linha2_3__48, linha2_3__47, linha2_3__46, linha2_3__45, 
         linha2_3__44, linha2_3__43, linha2_3__42, linha2_3__41, linha2_3__40, 
         linha2_3__39, linha2_3__38, linha2_3__37, linha2_3__36, linha2_3__35, 
         linha2_3__34, linha2_3__33, linha2_3__32, linha2_3__31, linha2_3__30, 
         linha2_3__29, linha2_3__28, linha2_3__27, linha2_3__26, linha2_3__25, 
         linha2_3__24, linha2_3__23, linha2_3__22, linha2_3__21, linha2_3__20, 
         linha2_3__19, linha2_3__18, linha2_3__17, linha2_3__16, linha2_3__15, 
         linha2_3__14, linha2_3__13, linha2_3__12, linha2_3__11, linha2_3__10, 
         linha2_3__9, linha2_3__8, linha2_3__7, linha2_3__6, linha2_3__5, 
         linha2_3__4, linha2_3__3, linha2_3__2, linha2_3__1, linha2_3__0, 
         linha2_2__63, linha2_2__62, linha2_2__61, linha2_2__60, linha2_2__59, 
         linha2_2__58, linha2_2__57, linha2_2__56, linha2_2__55, linha2_2__54, 
         linha2_2__53, linha2_2__52, linha2_2__51, linha2_2__50, linha2_2__49, 
         linha2_2__48, linha2_2__47, linha2_2__46, linha2_2__45, linha2_2__44, 
         linha2_2__43, linha2_2__42, linha2_2__41, linha2_2__40, linha2_2__39, 
         linha2_2__38, linha2_2__37, linha2_2__36, linha2_2__35, linha2_2__34, 
         linha2_2__33, linha2_2__32, linha2_2__31, linha2_2__30, linha2_2__29, 
         linha2_2__28, linha2_2__27, linha2_2__26, linha2_2__25, linha2_2__24, 
         linha2_2__23, linha2_2__22, linha2_2__21, linha2_2__20, linha2_2__19, 
         linha2_2__18, linha2_2__17, linha2_2__16, linha2_2__15, linha2_2__14, 
         linha2_2__13, linha2_2__12, linha2_2__11, linha2_2__10, linha2_2__9, 
         linha2_2__8, linha2_2__7, linha2_2__6, linha2_2__5, linha2_2__4, 
         linha2_2__3, linha2_2__2, linha2_2__1, linha2_2__0, linha2_1__63, 
         linha2_1__62, linha2_1__61, linha2_1__60, linha2_1__59, linha2_1__58, 
         linha2_1__57, linha2_1__56, linha2_1__55, linha2_1__54, linha2_1__53, 
         linha2_1__52, linha2_1__51, linha2_1__50, linha2_1__49, linha2_1__48, 
         linha2_1__47, linha2_1__46, linha2_1__45, linha2_1__44, linha2_1__43, 
         linha2_1__42, linha2_1__41, linha2_1__40, linha2_1__39, linha2_1__38, 
         linha2_1__37, linha2_1__36, linha2_1__35, linha2_1__34, linha2_1__33, 
         linha2_1__32, linha2_1__31, linha2_1__30, linha2_1__29, linha2_1__28, 
         linha2_1__27, linha2_1__26, linha2_1__25, linha2_1__24, linha2_1__23, 
         linha2_1__22, linha2_1__21, linha2_1__20, linha2_1__19, linha2_1__18, 
         linha2_1__17, linha2_1__16, linha2_1__15, linha2_1__14, linha2_1__13, 
         linha2_1__12, linha2_1__11, linha2_1__10, linha2_1__9, linha2_1__8, 
         linha2_1__7, linha2_1__6, linha2_1__5, linha2_1__4, linha2_1__3, 
         linha2_1__2, linha2_1__1, linha2_1__0, linha8_3__63, linha8_3__62, 
         linha8_3__61, linha8_3__60, linha8_3__59, linha8_3__58, linha8_3__57, 
         linha8_3__56, linha8_3__55, linha8_3__54, linha8_3__53, linha8_3__52, 
         linha8_3__51, linha8_3__50, linha8_3__49, linha8_3__48, linha8_3__47, 
         linha8_3__46, linha8_3__45, linha8_3__44, linha8_3__43, linha8_3__42, 
         linha8_3__41, linha8_3__40, linha8_3__39, linha8_3__38, linha8_3__37, 
         linha8_3__36, linha8_3__35, linha8_3__34, linha8_3__33, linha8_3__32, 
         linha8_3__31, linha8_3__30, linha8_3__29, linha8_3__28, linha8_3__27, 
         linha8_3__26, linha8_3__25, linha8_3__24, linha8_3__23, linha8_3__22, 
         linha8_3__21, linha8_3__20, linha8_3__19, linha8_3__18, linha8_3__17, 
         linha8_3__16, linha8_3__15, linha8_3__14, linha8_3__13, linha8_3__12, 
         linha8_3__11, linha8_3__10, linha8_3__9, linha8_3__8, linha8_3__7, 
         linha8_3__6, linha8_3__5, linha8_3__4, linha8_3__3, linha8_3__2, 
         linha8_3__1, linha8_3__0, linha8_2__63, linha8_2__62, linha8_2__61, 
         linha8_2__60, linha8_2__59, linha8_2__58, linha8_2__57, linha8_2__56, 
         linha8_2__55, linha8_2__54, linha8_2__53, linha8_2__52, linha8_2__51, 
         linha8_2__50, linha8_2__49, linha8_2__48, linha8_2__47, linha8_2__46, 
         linha8_2__45, linha8_2__44, linha8_2__43, linha8_2__42, linha8_2__41, 
         linha8_2__40, linha8_2__39, linha8_2__38, linha8_2__37, linha8_2__36, 
         linha8_2__35, linha8_2__34, linha8_2__33, linha8_2__32, linha8_2__31, 
         linha8_2__30, linha8_2__29, linha8_2__28, linha8_2__27, linha8_2__26, 
         linha8_2__25, linha8_2__24, linha8_2__23, linha8_2__22, linha8_2__21, 
         linha8_2__20, linha8_2__19, linha8_2__18, linha8_2__17, linha8_2__16, 
         linha8_2__15, linha8_2__14, linha8_2__13, linha8_2__12, linha8_2__11, 
         linha8_2__10, linha8_2__9, linha8_2__8, linha8_2__7, linha8_2__6, 
         linha8_2__5, linha8_2__4, linha8_2__3, linha8_2__2, linha8_2__1, 
         linha8_2__0, linha8_1__63, linha8_1__62, linha8_1__61, linha8_1__60, 
         linha8_1__59, linha8_1__58, linha8_1__57, linha8_1__56, linha8_1__55, 
         linha8_1__54, linha8_1__53, linha8_1__52, linha8_1__51, linha8_1__50, 
         linha8_1__49, linha8_1__48, linha8_1__47, linha8_1__46, linha8_1__45, 
         linha8_1__44, linha8_1__43, linha8_1__42, linha8_1__41, linha8_1__40, 
         linha8_1__39, linha8_1__38, linha8_1__37, linha8_1__36, linha8_1__35, 
         linha8_1__34, linha8_1__33, linha8_1__32, linha8_1__31, linha8_1__30, 
         linha8_1__29, linha8_1__28, linha8_1__27, linha8_1__26, linha8_1__25, 
         linha8_1__24, linha8_1__23, linha8_1__22, linha8_1__21, linha8_1__20, 
         linha8_1__19, linha8_1__18, linha8_1__17, linha8_1__16, linha8_1__15, 
         linha8_1__14, linha8_1__13, linha8_1__12, linha8_1__11, linha8_1__10, 
         linha8_1__9, linha8_1__8, linha8_1__7, linha8_1__6, linha8_1__5, 
         linha8_1__4, linha8_1__3, linha8_1__2, linha8_1__1, linha8_1__0, 
         linha1_3__63, linha1_3__62, linha1_3__61, linha1_3__60, linha1_3__59, 
         linha1_3__58, linha1_3__57, linha1_3__56, linha1_3__55, linha1_3__54, 
         linha1_3__53, linha1_3__52, linha1_3__51, linha1_3__50, linha1_3__49, 
         linha1_3__48, linha1_3__47, linha1_3__46, linha1_3__45, linha1_3__44, 
         linha1_3__43, linha1_3__42, linha1_3__41, linha1_3__40, linha1_3__39, 
         linha1_3__38, linha1_3__37, linha1_3__36, linha1_3__35, linha1_3__34, 
         linha1_3__33, linha1_3__32, linha1_3__31, linha1_3__30, linha1_3__29, 
         linha1_3__28, linha1_3__27, linha1_3__26, linha1_3__25, linha1_3__24, 
         linha1_3__23, linha1_3__22, linha1_3__21, linha1_3__20, linha1_3__19, 
         linha1_3__18, linha1_3__17, linha1_3__16, linha1_3__15, linha1_3__14, 
         linha1_3__13, linha1_3__12, linha1_3__11, linha1_3__10, linha1_3__9, 
         linha1_3__8, linha1_3__7, linha1_3__6, linha1_3__5, linha1_3__4, 
         linha1_3__3, linha1_3__2, linha1_3__1, linha1_3__0, linha1_2__63, 
         linha1_2__62, linha1_2__61, linha1_2__60, linha1_2__59, linha1_2__58, 
         linha1_2__57, linha1_2__56, linha1_2__55, linha1_2__54, linha1_2__53, 
         linha1_2__52, linha1_2__51, linha1_2__50, linha1_2__49, linha1_2__48, 
         linha1_2__47, linha1_2__46, linha1_2__45, linha1_2__44, linha1_2__43, 
         linha1_2__42, linha1_2__41, linha1_2__40, linha1_2__39, linha1_2__38, 
         linha1_2__37, linha1_2__36, linha1_2__35, linha1_2__34, linha1_2__33, 
         linha1_2__32, linha1_2__31, linha1_2__30, linha1_2__29, linha1_2__28, 
         linha1_2__27, linha1_2__26, linha1_2__25, linha1_2__24, linha1_2__23, 
         linha1_2__22, linha1_2__21, linha1_2__20, linha1_2__19, linha1_2__18, 
         linha1_2__17, linha1_2__16, linha1_2__15, linha1_2__14, linha1_2__13, 
         linha1_2__12, linha1_2__11, linha1_2__10, linha1_2__9, linha1_2__8, 
         linha1_2__7, linha1_2__6, linha1_2__5, linha1_2__4, linha1_2__3, 
         linha1_2__2, linha1_2__1, linha1_2__0, linha1_1__63, linha1_1__62, 
         linha1_1__61, linha1_1__60, linha1_1__59, linha1_1__58, linha1_1__57, 
         linha1_1__56, linha1_1__55, linha1_1__54, linha1_1__53, linha1_1__52, 
         linha1_1__51, linha1_1__50, linha1_1__49, linha1_1__48, linha1_1__47, 
         linha1_1__46, linha1_1__45, linha1_1__44, linha1_1__43, linha1_1__42, 
         linha1_1__41, linha1_1__40, linha1_1__39, linha1_1__38, linha1_1__37, 
         linha1_1__36, linha1_1__35, linha1_1__34, linha1_1__33, linha1_1__32, 
         linha1_1__31, linha1_1__30, linha1_1__29, linha1_1__28, linha1_1__27, 
         linha1_1__26, linha1_1__25, linha1_1__24, linha1_1__23, linha1_1__22, 
         linha1_1__21, linha1_1__20, linha1_1__19, linha1_1__18, linha1_1__17, 
         linha1_1__16, linha1_1__15, linha1_1__14, linha1_1__13, linha1_1__12, 
         linha1_1__11, linha1_1__10, linha1_1__9, linha1_1__8, linha1_1__7, 
         linha1_1__6, linha1_1__5, linha1_1__4, linha1_1__3, linha1_1__2, 
         linha1_1__1, linha1_1__0, row_0_rowp_bni1_l, row_0_rowp_bni2_l, 
         row_0_rowp_bni3_l, row_0_rowp_bni4_l, row_1_rowi_bni1_l, 
         row_1_rowi_bni2_l, row_1_rowi_bni3_l, row_2_rowp_bni1_l, 
         row_2_rowp_bni2_l, row_2_rowp_bni3_l, row_2_rowp_bni4_l, 
         row_3_rowi_bni1_l, row_3_rowi_bni2_l, row_3_rowi_bni3_l, 
         row_4_rowp_bni1_l, row_4_rowp_bni2_l, row_4_rowp_bni3_l, 
         row_4_rowp_bni4_l, row_5_rowi_bni1_l, row_5_rowi_bni2_l, 
         row_5_rowi_bni3_l, row_6_rowp_bni1_l, row_6_rowp_bni2_l, 
         row_6_rowp_bni3_l, row_6_rowp_bni4_l, row_7_rowi_bni1_l, 
         row_7_rowi_bni2_l, row_7_rowi_bni3_l, nx8127;
    wire [27:0] \$dummy ;




    juntarComparadores_64 row_0_rowp_bni1_Comp (.g (\$dummy [0]), .l (
                          row_0_rowp_bni1_l), .a ({x1[63],x1[62],x1[61],x1[60],
                          x1[59],x1[58],x1[57],x1[56],x1[55],x1[54],x1[53],
                          x1[52],x1[51],x1[50],x1[49],x1[48],x1[47],x1[46],
                          x1[45],x1[44],x1[43],x1[42],x1[41],x1[40],x1[39],
                          x1[38],x1[37],x1[36],x1[35],x1[34],x1[33],x1[32],
                          x1[31],x1[30],x1[29],x1[28],x1[27],x1[26],x1[25],
                          x1[24],x1[23],x1[22],x1[21],x1[20],x1[19],x1[18],
                          x1[17],x1[16],x1[15],x1[14],x1[13],x1[12],x1[11],
                          x1[10],x1[9],x1[8],x1[7],x1[6],x1[5],x1[4],x1[3],x1[2]
                          ,x1[1],x1[0]}), .b ({x2[63],x2[62],x2[61],x2[60],
                          x2[59],x2[58],x2[57],x2[56],x2[55],x2[54],x2[53],
                          x2[52],x2[51],x2[50],x2[49],x2[48],x2[47],x2[46],
                          x2[45],x2[44],x2[43],x2[42],x2[41],x2[40],x2[39],
                          x2[38],x2[37],x2[36],x2[35],x2[34],x2[33],x2[32],
                          x2[31],x2[30],x2[29],x2[28],x2[27],x2[26],x2[25],
                          x2[24],x2[23],x2[22],x2[21],x2[20],x2[19],x2[18],
                          x2[17],x2[16],x2[15],x2[14],x2[13],x2[12],x2[11],
                          x2[10],x2[9],x2[8],x2[7],x2[6],x2[5],x2[4],x2[3],x2[2]
                          ,x2[1],x2[0]})) ;
    Mux2x1_64 row_0_rowp_bni1_muxMax (.r ({linha1_1__63,linha1_1__62,
              linha1_1__61,linha1_1__60,linha1_1__59,linha1_1__58,linha1_1__57,
              linha1_1__56,linha1_1__55,linha1_1__54,linha1_1__53,linha1_1__52,
              linha1_1__51,linha1_1__50,linha1_1__49,linha1_1__48,linha1_1__47,
              linha1_1__46,linha1_1__45,linha1_1__44,linha1_1__43,linha1_1__42,
              linha1_1__41,linha1_1__40,linha1_1__39,linha1_1__38,linha1_1__37,
              linha1_1__36,linha1_1__35,linha1_1__34,linha1_1__33,linha1_1__32,
              linha1_1__31,linha1_1__30,linha1_1__29,linha1_1__28,linha1_1__27,
              linha1_1__26,linha1_1__25,linha1_1__24,linha1_1__23,linha1_1__22,
              linha1_1__21,linha1_1__20,linha1_1__19,linha1_1__18,linha1_1__17,
              linha1_1__16,linha1_1__15,linha1_1__14,linha1_1__13,linha1_1__12,
              linha1_1__11,linha1_1__10,linha1_1__9,linha1_1__8,linha1_1__7,
              linha1_1__6,linha1_1__5,linha1_1__4,linha1_1__3,linha1_1__2,
              linha1_1__1,linha1_1__0}), .a1 ({x2[63],x2[62],x2[61],x2[60],
              x2[59],x2[58],x2[57],x2[56],x2[55],x2[54],x2[53],x2[52],x2[51],
              x2[50],x2[49],x2[48],x2[47],x2[46],x2[45],x2[44],x2[43],x2[42],
              x2[41],x2[40],x2[39],x2[38],x2[37],x2[36],x2[35],x2[34],x2[33],
              x2[32],x2[31],x2[30],x2[29],x2[28],x2[27],x2[26],x2[25],x2[24],
              x2[23],x2[22],x2[21],x2[20],x2[19],x2[18],x2[17],x2[16],x2[15],
              x2[14],x2[13],x2[12],x2[11],x2[10],x2[9],x2[8],x2[7],x2[6],x2[5],
              x2[4],x2[3],x2[2],x2[1],x2[0]}), .a0 ({x1[63],x1[62],x1[61],x1[60]
              ,x1[59],x1[58],x1[57],x1[56],x1[55],x1[54],x1[53],x1[52],x1[51],
              x1[50],x1[49],x1[48],x1[47],x1[46],x1[45],x1[44],x1[43],x1[42],
              x1[41],x1[40],x1[39],x1[38],x1[37],x1[36],x1[35],x1[34],x1[33],
              x1[32],x1[31],x1[30],x1[29],x1[28],x1[27],x1[26],x1[25],x1[24],
              x1[23],x1[22],x1[21],x1[20],x1[19],x1[18],x1[17],x1[16],x1[15],
              x1[14],x1[13],x1[12],x1[11],x1[10],x1[9],x1[8],x1[7],x1[6],x1[5],
              x1[4],x1[3],x1[2],x1[1],x1[0]}), .s (nx8127)) ;
    Mux2x1_64 row_0_rowp_bni1_muxMin (.r ({linha2_1__63,linha2_1__62,
              linha2_1__61,linha2_1__60,linha2_1__59,linha2_1__58,linha2_1__57,
              linha2_1__56,linha2_1__55,linha2_1__54,linha2_1__53,linha2_1__52,
              linha2_1__51,linha2_1__50,linha2_1__49,linha2_1__48,linha2_1__47,
              linha2_1__46,linha2_1__45,linha2_1__44,linha2_1__43,linha2_1__42,
              linha2_1__41,linha2_1__40,linha2_1__39,linha2_1__38,linha2_1__37,
              linha2_1__36,linha2_1__35,linha2_1__34,linha2_1__33,linha2_1__32,
              linha2_1__31,linha2_1__30,linha2_1__29,linha2_1__28,linha2_1__27,
              linha2_1__26,linha2_1__25,linha2_1__24,linha2_1__23,linha2_1__22,
              linha2_1__21,linha2_1__20,linha2_1__19,linha2_1__18,linha2_1__17,
              linha2_1__16,linha2_1__15,linha2_1__14,linha2_1__13,linha2_1__12,
              linha2_1__11,linha2_1__10,linha2_1__9,linha2_1__8,linha2_1__7,
              linha2_1__6,linha2_1__5,linha2_1__4,linha2_1__3,linha2_1__2,
              linha2_1__1,linha2_1__0}), .a1 ({x1[63],x1[62],x1[61],x1[60],
              x1[59],x1[58],x1[57],x1[56],x1[55],x1[54],x1[53],x1[52],x1[51],
              x1[50],x1[49],x1[48],x1[47],x1[46],x1[45],x1[44],x1[43],x1[42],
              x1[41],x1[40],x1[39],x1[38],x1[37],x1[36],x1[35],x1[34],x1[33],
              x1[32],x1[31],x1[30],x1[29],x1[28],x1[27],x1[26],x1[25],x1[24],
              x1[23],x1[22],x1[21],x1[20],x1[19],x1[18],x1[17],x1[16],x1[15],
              x1[14],x1[13],x1[12],x1[11],x1[10],x1[9],x1[8],x1[7],x1[6],x1[5],
              x1[4],x1[3],x1[2],x1[1],x1[0]}), .a0 ({x2[63],x2[62],x2[61],x2[60]
              ,x2[59],x2[58],x2[57],x2[56],x2[55],x2[54],x2[53],x2[52],x2[51],
              x2[50],x2[49],x2[48],x2[47],x2[46],x2[45],x2[44],x2[43],x2[42],
              x2[41],x2[40],x2[39],x2[38],x2[37],x2[36],x2[35],x2[34],x2[33],
              x2[32],x2[31],x2[30],x2[29],x2[28],x2[27],x2[26],x2[25],x2[24],
              x2[23],x2[22],x2[21],x2[20],x2[19],x2[18],x2[17],x2[16],x2[15],
              x2[14],x2[13],x2[12],x2[11],x2[10],x2[9],x2[8],x2[7],x2[6],x2[5],
              x2[4],x2[3],x2[2],x2[1],x2[0]}), .s (nx8127)) ;
    juntarComparadores_64 row_0_rowp_bni2_Comp (.g (\$dummy [1]), .l (
                          row_0_rowp_bni2_l), .a ({x3[63],x3[62],x3[61],x3[60],
                          x3[59],x3[58],x3[57],x3[56],x3[55],x3[54],x3[53],
                          x3[52],x3[51],x3[50],x3[49],x3[48],x3[47],x3[46],
                          x3[45],x3[44],x3[43],x3[42],x3[41],x3[40],x3[39],
                          x3[38],x3[37],x3[36],x3[35],x3[34],x3[33],x3[32],
                          x3[31],x3[30],x3[29],x3[28],x3[27],x3[26],x3[25],
                          x3[24],x3[23],x3[22],x3[21],x3[20],x3[19],x3[18],
                          x3[17],x3[16],x3[15],x3[14],x3[13],x3[12],x3[11],
                          x3[10],x3[9],x3[8],x3[7],x3[6],x3[5],x3[4],x3[3],x3[2]
                          ,x3[1],x3[0]}), .b ({x4[63],x4[62],x4[61],x4[60],
                          x4[59],x4[58],x4[57],x4[56],x4[55],x4[54],x4[53],
                          x4[52],x4[51],x4[50],x4[49],x4[48],x4[47],x4[46],
                          x4[45],x4[44],x4[43],x4[42],x4[41],x4[40],x4[39],
                          x4[38],x4[37],x4[36],x4[35],x4[34],x4[33],x4[32],
                          x4[31],x4[30],x4[29],x4[28],x4[27],x4[26],x4[25],
                          x4[24],x4[23],x4[22],x4[21],x4[20],x4[19],x4[18],
                          x4[17],x4[16],x4[15],x4[14],x4[13],x4[12],x4[11],
                          x4[10],x4[9],x4[8],x4[7],x4[6],x4[5],x4[4],x4[3],x4[2]
                          ,x4[1],x4[0]})) ;
    Mux2x1_64 row_0_rowp_bni2_muxMax (.r ({linha3_1__63,linha3_1__62,
              linha3_1__61,linha3_1__60,linha3_1__59,linha3_1__58,linha3_1__57,
              linha3_1__56,linha3_1__55,linha3_1__54,linha3_1__53,linha3_1__52,
              linha3_1__51,linha3_1__50,linha3_1__49,linha3_1__48,linha3_1__47,
              linha3_1__46,linha3_1__45,linha3_1__44,linha3_1__43,linha3_1__42,
              linha3_1__41,linha3_1__40,linha3_1__39,linha3_1__38,linha3_1__37,
              linha3_1__36,linha3_1__35,linha3_1__34,linha3_1__33,linha3_1__32,
              linha3_1__31,linha3_1__30,linha3_1__29,linha3_1__28,linha3_1__27,
              linha3_1__26,linha3_1__25,linha3_1__24,linha3_1__23,linha3_1__22,
              linha3_1__21,linha3_1__20,linha3_1__19,linha3_1__18,linha3_1__17,
              linha3_1__16,linha3_1__15,linha3_1__14,linha3_1__13,linha3_1__12,
              linha3_1__11,linha3_1__10,linha3_1__9,linha3_1__8,linha3_1__7,
              linha3_1__6,linha3_1__5,linha3_1__4,linha3_1__3,linha3_1__2,
              linha3_1__1,linha3_1__0}), .a1 ({x4[63],x4[62],x4[61],x4[60],
              x4[59],x4[58],x4[57],x4[56],x4[55],x4[54],x4[53],x4[52],x4[51],
              x4[50],x4[49],x4[48],x4[47],x4[46],x4[45],x4[44],x4[43],x4[42],
              x4[41],x4[40],x4[39],x4[38],x4[37],x4[36],x4[35],x4[34],x4[33],
              x4[32],x4[31],x4[30],x4[29],x4[28],x4[27],x4[26],x4[25],x4[24],
              x4[23],x4[22],x4[21],x4[20],x4[19],x4[18],x4[17],x4[16],x4[15],
              x4[14],x4[13],x4[12],x4[11],x4[10],x4[9],x4[8],x4[7],x4[6],x4[5],
              x4[4],x4[3],x4[2],x4[1],x4[0]}), .a0 ({x3[63],x3[62],x3[61],x3[60]
              ,x3[59],x3[58],x3[57],x3[56],x3[55],x3[54],x3[53],x3[52],x3[51],
              x3[50],x3[49],x3[48],x3[47],x3[46],x3[45],x3[44],x3[43],x3[42],
              x3[41],x3[40],x3[39],x3[38],x3[37],x3[36],x3[35],x3[34],x3[33],
              x3[32],x3[31],x3[30],x3[29],x3[28],x3[27],x3[26],x3[25],x3[24],
              x3[23],x3[22],x3[21],x3[20],x3[19],x3[18],x3[17],x3[16],x3[15],
              x3[14],x3[13],x3[12],x3[11],x3[10],x3[9],x3[8],x3[7],x3[6],x3[5],
              x3[4],x3[3],x3[2],x3[1],x3[0]}), .s (row_0_rowp_bni2_l)) ;
    Mux2x1_64 row_0_rowp_bni2_muxMin (.r ({linha4_1__63,linha4_1__62,
              linha4_1__61,linha4_1__60,linha4_1__59,linha4_1__58,linha4_1__57,
              linha4_1__56,linha4_1__55,linha4_1__54,linha4_1__53,linha4_1__52,
              linha4_1__51,linha4_1__50,linha4_1__49,linha4_1__48,linha4_1__47,
              linha4_1__46,linha4_1__45,linha4_1__44,linha4_1__43,linha4_1__42,
              linha4_1__41,linha4_1__40,linha4_1__39,linha4_1__38,linha4_1__37,
              linha4_1__36,linha4_1__35,linha4_1__34,linha4_1__33,linha4_1__32,
              linha4_1__31,linha4_1__30,linha4_1__29,linha4_1__28,linha4_1__27,
              linha4_1__26,linha4_1__25,linha4_1__24,linha4_1__23,linha4_1__22,
              linha4_1__21,linha4_1__20,linha4_1__19,linha4_1__18,linha4_1__17,
              linha4_1__16,linha4_1__15,linha4_1__14,linha4_1__13,linha4_1__12,
              linha4_1__11,linha4_1__10,linha4_1__9,linha4_1__8,linha4_1__7,
              linha4_1__6,linha4_1__5,linha4_1__4,linha4_1__3,linha4_1__2,
              linha4_1__1,linha4_1__0}), .a1 ({x3[63],x3[62],x3[61],x3[60],
              x3[59],x3[58],x3[57],x3[56],x3[55],x3[54],x3[53],x3[52],x3[51],
              x3[50],x3[49],x3[48],x3[47],x3[46],x3[45],x3[44],x3[43],x3[42],
              x3[41],x3[40],x3[39],x3[38],x3[37],x3[36],x3[35],x3[34],x3[33],
              x3[32],x3[31],x3[30],x3[29],x3[28],x3[27],x3[26],x3[25],x3[24],
              x3[23],x3[22],x3[21],x3[20],x3[19],x3[18],x3[17],x3[16],x3[15],
              x3[14],x3[13],x3[12],x3[11],x3[10],x3[9],x3[8],x3[7],x3[6],x3[5],
              x3[4],x3[3],x3[2],x3[1],x3[0]}), .a0 ({x4[63],x4[62],x4[61],x4[60]
              ,x4[59],x4[58],x4[57],x4[56],x4[55],x4[54],x4[53],x4[52],x4[51],
              x4[50],x4[49],x4[48],x4[47],x4[46],x4[45],x4[44],x4[43],x4[42],
              x4[41],x4[40],x4[39],x4[38],x4[37],x4[36],x4[35],x4[34],x4[33],
              x4[32],x4[31],x4[30],x4[29],x4[28],x4[27],x4[26],x4[25],x4[24],
              x4[23],x4[22],x4[21],x4[20],x4[19],x4[18],x4[17],x4[16],x4[15],
              x4[14],x4[13],x4[12],x4[11],x4[10],x4[9],x4[8],x4[7],x4[6],x4[5],
              x4[4],x4[3],x4[2],x4[1],x4[0]}), .s (row_0_rowp_bni2_l)) ;
    juntarComparadores_64 row_0_rowp_bni3_Comp (.g (\$dummy [2]), .l (
                          row_0_rowp_bni3_l), .a ({x5[63],x5[62],x5[61],x5[60],
                          x5[59],x5[58],x5[57],x5[56],x5[55],x5[54],x5[53],
                          x5[52],x5[51],x5[50],x5[49],x5[48],x5[47],x5[46],
                          x5[45],x5[44],x5[43],x5[42],x5[41],x5[40],x5[39],
                          x5[38],x5[37],x5[36],x5[35],x5[34],x5[33],x5[32],
                          x5[31],x5[30],x5[29],x5[28],x5[27],x5[26],x5[25],
                          x5[24],x5[23],x5[22],x5[21],x5[20],x5[19],x5[18],
                          x5[17],x5[16],x5[15],x5[14],x5[13],x5[12],x5[11],
                          x5[10],x5[9],x5[8],x5[7],x5[6],x5[5],x5[4],x5[3],x5[2]
                          ,x5[1],x5[0]}), .b ({x6[63],x6[62],x6[61],x6[60],
                          x6[59],x6[58],x6[57],x6[56],x6[55],x6[54],x6[53],
                          x6[52],x6[51],x6[50],x6[49],x6[48],x6[47],x6[46],
                          x6[45],x6[44],x6[43],x6[42],x6[41],x6[40],x6[39],
                          x6[38],x6[37],x6[36],x6[35],x6[34],x6[33],x6[32],
                          x6[31],x6[30],x6[29],x6[28],x6[27],x6[26],x6[25],
                          x6[24],x6[23],x6[22],x6[21],x6[20],x6[19],x6[18],
                          x6[17],x6[16],x6[15],x6[14],x6[13],x6[12],x6[11],
                          x6[10],x6[9],x6[8],x6[7],x6[6],x6[5],x6[4],x6[3],x6[2]
                          ,x6[1],x6[0]})) ;
    Mux2x1_64 row_0_rowp_bni3_muxMax (.r ({linha5_1__63,linha5_1__62,
              linha5_1__61,linha5_1__60,linha5_1__59,linha5_1__58,linha5_1__57,
              linha5_1__56,linha5_1__55,linha5_1__54,linha5_1__53,linha5_1__52,
              linha5_1__51,linha5_1__50,linha5_1__49,linha5_1__48,linha5_1__47,
              linha5_1__46,linha5_1__45,linha5_1__44,linha5_1__43,linha5_1__42,
              linha5_1__41,linha5_1__40,linha5_1__39,linha5_1__38,linha5_1__37,
              linha5_1__36,linha5_1__35,linha5_1__34,linha5_1__33,linha5_1__32,
              linha5_1__31,linha5_1__30,linha5_1__29,linha5_1__28,linha5_1__27,
              linha5_1__26,linha5_1__25,linha5_1__24,linha5_1__23,linha5_1__22,
              linha5_1__21,linha5_1__20,linha5_1__19,linha5_1__18,linha5_1__17,
              linha5_1__16,linha5_1__15,linha5_1__14,linha5_1__13,linha5_1__12,
              linha5_1__11,linha5_1__10,linha5_1__9,linha5_1__8,linha5_1__7,
              linha5_1__6,linha5_1__5,linha5_1__4,linha5_1__3,linha5_1__2,
              linha5_1__1,linha5_1__0}), .a1 ({x6[63],x6[62],x6[61],x6[60],
              x6[59],x6[58],x6[57],x6[56],x6[55],x6[54],x6[53],x6[52],x6[51],
              x6[50],x6[49],x6[48],x6[47],x6[46],x6[45],x6[44],x6[43],x6[42],
              x6[41],x6[40],x6[39],x6[38],x6[37],x6[36],x6[35],x6[34],x6[33],
              x6[32],x6[31],x6[30],x6[29],x6[28],x6[27],x6[26],x6[25],x6[24],
              x6[23],x6[22],x6[21],x6[20],x6[19],x6[18],x6[17],x6[16],x6[15],
              x6[14],x6[13],x6[12],x6[11],x6[10],x6[9],x6[8],x6[7],x6[6],x6[5],
              x6[4],x6[3],x6[2],x6[1],x6[0]}), .a0 ({x5[63],x5[62],x5[61],x5[60]
              ,x5[59],x5[58],x5[57],x5[56],x5[55],x5[54],x5[53],x5[52],x5[51],
              x5[50],x5[49],x5[48],x5[47],x5[46],x5[45],x5[44],x5[43],x5[42],
              x5[41],x5[40],x5[39],x5[38],x5[37],x5[36],x5[35],x5[34],x5[33],
              x5[32],x5[31],x5[30],x5[29],x5[28],x5[27],x5[26],x5[25],x5[24],
              x5[23],x5[22],x5[21],x5[20],x5[19],x5[18],x5[17],x5[16],x5[15],
              x5[14],x5[13],x5[12],x5[11],x5[10],x5[9],x5[8],x5[7],x5[6],x5[5],
              x5[4],x5[3],x5[2],x5[1],x5[0]}), .s (row_0_rowp_bni3_l)) ;
    Mux2x1_64 row_0_rowp_bni3_muxMin (.r ({linha6_1__63,linha6_1__62,
              linha6_1__61,linha6_1__60,linha6_1__59,linha6_1__58,linha6_1__57,
              linha6_1__56,linha6_1__55,linha6_1__54,linha6_1__53,linha6_1__52,
              linha6_1__51,linha6_1__50,linha6_1__49,linha6_1__48,linha6_1__47,
              linha6_1__46,linha6_1__45,linha6_1__44,linha6_1__43,linha6_1__42,
              linha6_1__41,linha6_1__40,linha6_1__39,linha6_1__38,linha6_1__37,
              linha6_1__36,linha6_1__35,linha6_1__34,linha6_1__33,linha6_1__32,
              linha6_1__31,linha6_1__30,linha6_1__29,linha6_1__28,linha6_1__27,
              linha6_1__26,linha6_1__25,linha6_1__24,linha6_1__23,linha6_1__22,
              linha6_1__21,linha6_1__20,linha6_1__19,linha6_1__18,linha6_1__17,
              linha6_1__16,linha6_1__15,linha6_1__14,linha6_1__13,linha6_1__12,
              linha6_1__11,linha6_1__10,linha6_1__9,linha6_1__8,linha6_1__7,
              linha6_1__6,linha6_1__5,linha6_1__4,linha6_1__3,linha6_1__2,
              linha6_1__1,linha6_1__0}), .a1 ({x5[63],x5[62],x5[61],x5[60],
              x5[59],x5[58],x5[57],x5[56],x5[55],x5[54],x5[53],x5[52],x5[51],
              x5[50],x5[49],x5[48],x5[47],x5[46],x5[45],x5[44],x5[43],x5[42],
              x5[41],x5[40],x5[39],x5[38],x5[37],x5[36],x5[35],x5[34],x5[33],
              x5[32],x5[31],x5[30],x5[29],x5[28],x5[27],x5[26],x5[25],x5[24],
              x5[23],x5[22],x5[21],x5[20],x5[19],x5[18],x5[17],x5[16],x5[15],
              x5[14],x5[13],x5[12],x5[11],x5[10],x5[9],x5[8],x5[7],x5[6],x5[5],
              x5[4],x5[3],x5[2],x5[1],x5[0]}), .a0 ({x6[63],x6[62],x6[61],x6[60]
              ,x6[59],x6[58],x6[57],x6[56],x6[55],x6[54],x6[53],x6[52],x6[51],
              x6[50],x6[49],x6[48],x6[47],x6[46],x6[45],x6[44],x6[43],x6[42],
              x6[41],x6[40],x6[39],x6[38],x6[37],x6[36],x6[35],x6[34],x6[33],
              x6[32],x6[31],x6[30],x6[29],x6[28],x6[27],x6[26],x6[25],x6[24],
              x6[23],x6[22],x6[21],x6[20],x6[19],x6[18],x6[17],x6[16],x6[15],
              x6[14],x6[13],x6[12],x6[11],x6[10],x6[9],x6[8],x6[7],x6[6],x6[5],
              x6[4],x6[3],x6[2],x6[1],x6[0]}), .s (row_0_rowp_bni3_l)) ;
    juntarComparadores_64 row_0_rowp_bni4_Comp (.g (\$dummy [3]), .l (
                          row_0_rowp_bni4_l), .a ({x7[63],x7[62],x7[61],x7[60],
                          x7[59],x7[58],x7[57],x7[56],x7[55],x7[54],x7[53],
                          x7[52],x7[51],x7[50],x7[49],x7[48],x7[47],x7[46],
                          x7[45],x7[44],x7[43],x7[42],x7[41],x7[40],x7[39],
                          x7[38],x7[37],x7[36],x7[35],x7[34],x7[33],x7[32],
                          x7[31],x7[30],x7[29],x7[28],x7[27],x7[26],x7[25],
                          x7[24],x7[23],x7[22],x7[21],x7[20],x7[19],x7[18],
                          x7[17],x7[16],x7[15],x7[14],x7[13],x7[12],x7[11],
                          x7[10],x7[9],x7[8],x7[7],x7[6],x7[5],x7[4],x7[3],x7[2]
                          ,x7[1],x7[0]}), .b ({x8[63],x8[62],x8[61],x8[60],
                          x8[59],x8[58],x8[57],x8[56],x8[55],x8[54],x8[53],
                          x8[52],x8[51],x8[50],x8[49],x8[48],x8[47],x8[46],
                          x8[45],x8[44],x8[43],x8[42],x8[41],x8[40],x8[39],
                          x8[38],x8[37],x8[36],x8[35],x8[34],x8[33],x8[32],
                          x8[31],x8[30],x8[29],x8[28],x8[27],x8[26],x8[25],
                          x8[24],x8[23],x8[22],x8[21],x8[20],x8[19],x8[18],
                          x8[17],x8[16],x8[15],x8[14],x8[13],x8[12],x8[11],
                          x8[10],x8[9],x8[8],x8[7],x8[6],x8[5],x8[4],x8[3],x8[2]
                          ,x8[1],x8[0]})) ;
    Mux2x1_64 row_0_rowp_bni4_muxMax (.r ({linha7_1__63,linha7_1__62,
              linha7_1__61,linha7_1__60,linha7_1__59,linha7_1__58,linha7_1__57,
              linha7_1__56,linha7_1__55,linha7_1__54,linha7_1__53,linha7_1__52,
              linha7_1__51,linha7_1__50,linha7_1__49,linha7_1__48,linha7_1__47,
              linha7_1__46,linha7_1__45,linha7_1__44,linha7_1__43,linha7_1__42,
              linha7_1__41,linha7_1__40,linha7_1__39,linha7_1__38,linha7_1__37,
              linha7_1__36,linha7_1__35,linha7_1__34,linha7_1__33,linha7_1__32,
              linha7_1__31,linha7_1__30,linha7_1__29,linha7_1__28,linha7_1__27,
              linha7_1__26,linha7_1__25,linha7_1__24,linha7_1__23,linha7_1__22,
              linha7_1__21,linha7_1__20,linha7_1__19,linha7_1__18,linha7_1__17,
              linha7_1__16,linha7_1__15,linha7_1__14,linha7_1__13,linha7_1__12,
              linha7_1__11,linha7_1__10,linha7_1__9,linha7_1__8,linha7_1__7,
              linha7_1__6,linha7_1__5,linha7_1__4,linha7_1__3,linha7_1__2,
              linha7_1__1,linha7_1__0}), .a1 ({x8[63],x8[62],x8[61],x8[60],
              x8[59],x8[58],x8[57],x8[56],x8[55],x8[54],x8[53],x8[52],x8[51],
              x8[50],x8[49],x8[48],x8[47],x8[46],x8[45],x8[44],x8[43],x8[42],
              x8[41],x8[40],x8[39],x8[38],x8[37],x8[36],x8[35],x8[34],x8[33],
              x8[32],x8[31],x8[30],x8[29],x8[28],x8[27],x8[26],x8[25],x8[24],
              x8[23],x8[22],x8[21],x8[20],x8[19],x8[18],x8[17],x8[16],x8[15],
              x8[14],x8[13],x8[12],x8[11],x8[10],x8[9],x8[8],x8[7],x8[6],x8[5],
              x8[4],x8[3],x8[2],x8[1],x8[0]}), .a0 ({x7[63],x7[62],x7[61],x7[60]
              ,x7[59],x7[58],x7[57],x7[56],x7[55],x7[54],x7[53],x7[52],x7[51],
              x7[50],x7[49],x7[48],x7[47],x7[46],x7[45],x7[44],x7[43],x7[42],
              x7[41],x7[40],x7[39],x7[38],x7[37],x7[36],x7[35],x7[34],x7[33],
              x7[32],x7[31],x7[30],x7[29],x7[28],x7[27],x7[26],x7[25],x7[24],
              x7[23],x7[22],x7[21],x7[20],x7[19],x7[18],x7[17],x7[16],x7[15],
              x7[14],x7[13],x7[12],x7[11],x7[10],x7[9],x7[8],x7[7],x7[6],x7[5],
              x7[4],x7[3],x7[2],x7[1],x7[0]}), .s (row_0_rowp_bni4_l)) ;
    Mux2x1_64 row_0_rowp_bni4_muxMin (.r ({linha8_1__63,linha8_1__62,
              linha8_1__61,linha8_1__60,linha8_1__59,linha8_1__58,linha8_1__57,
              linha8_1__56,linha8_1__55,linha8_1__54,linha8_1__53,linha8_1__52,
              linha8_1__51,linha8_1__50,linha8_1__49,linha8_1__48,linha8_1__47,
              linha8_1__46,linha8_1__45,linha8_1__44,linha8_1__43,linha8_1__42,
              linha8_1__41,linha8_1__40,linha8_1__39,linha8_1__38,linha8_1__37,
              linha8_1__36,linha8_1__35,linha8_1__34,linha8_1__33,linha8_1__32,
              linha8_1__31,linha8_1__30,linha8_1__29,linha8_1__28,linha8_1__27,
              linha8_1__26,linha8_1__25,linha8_1__24,linha8_1__23,linha8_1__22,
              linha8_1__21,linha8_1__20,linha8_1__19,linha8_1__18,linha8_1__17,
              linha8_1__16,linha8_1__15,linha8_1__14,linha8_1__13,linha8_1__12,
              linha8_1__11,linha8_1__10,linha8_1__9,linha8_1__8,linha8_1__7,
              linha8_1__6,linha8_1__5,linha8_1__4,linha8_1__3,linha8_1__2,
              linha8_1__1,linha8_1__0}), .a1 ({x7[63],x7[62],x7[61],x7[60],
              x7[59],x7[58],x7[57],x7[56],x7[55],x7[54],x7[53],x7[52],x7[51],
              x7[50],x7[49],x7[48],x7[47],x7[46],x7[45],x7[44],x7[43],x7[42],
              x7[41],x7[40],x7[39],x7[38],x7[37],x7[36],x7[35],x7[34],x7[33],
              x7[32],x7[31],x7[30],x7[29],x7[28],x7[27],x7[26],x7[25],x7[24],
              x7[23],x7[22],x7[21],x7[20],x7[19],x7[18],x7[17],x7[16],x7[15],
              x7[14],x7[13],x7[12],x7[11],x7[10],x7[9],x7[8],x7[7],x7[6],x7[5],
              x7[4],x7[3],x7[2],x7[1],x7[0]}), .a0 ({x8[63],x8[62],x8[61],x8[60]
              ,x8[59],x8[58],x8[57],x8[56],x8[55],x8[54],x8[53],x8[52],x8[51],
              x8[50],x8[49],x8[48],x8[47],x8[46],x8[45],x8[44],x8[43],x8[42],
              x8[41],x8[40],x8[39],x8[38],x8[37],x8[36],x8[35],x8[34],x8[33],
              x8[32],x8[31],x8[30],x8[29],x8[28],x8[27],x8[26],x8[25],x8[24],
              x8[23],x8[22],x8[21],x8[20],x8[19],x8[18],x8[17],x8[16],x8[15],
              x8[14],x8[13],x8[12],x8[11],x8[10],x8[9],x8[8],x8[7],x8[6],x8[5],
              x8[4],x8[3],x8[2],x8[1],x8[0]}), .s (row_0_rowp_bni4_l)) ;
    juntarComparadores_64 row_1_rowi_bni1_Comp (.g (\$dummy [4]), .l (
                          row_1_rowi_bni1_l), .a ({linha2_1__63,linha2_1__62,
                          linha2_1__61,linha2_1__60,linha2_1__59,linha2_1__58,
                          linha2_1__57,linha2_1__56,linha2_1__55,linha2_1__54,
                          linha2_1__53,linha2_1__52,linha2_1__51,linha2_1__50,
                          linha2_1__49,linha2_1__48,linha2_1__47,linha2_1__46,
                          linha2_1__45,linha2_1__44,linha2_1__43,linha2_1__42,
                          linha2_1__41,linha2_1__40,linha2_1__39,linha2_1__38,
                          linha2_1__37,linha2_1__36,linha2_1__35,linha2_1__34,
                          linha2_1__33,linha2_1__32,linha2_1__31,linha2_1__30,
                          linha2_1__29,linha2_1__28,linha2_1__27,linha2_1__26,
                          linha2_1__25,linha2_1__24,linha2_1__23,linha2_1__22,
                          linha2_1__21,linha2_1__20,linha2_1__19,linha2_1__18,
                          linha2_1__17,linha2_1__16,linha2_1__15,linha2_1__14,
                          linha2_1__13,linha2_1__12,linha2_1__11,linha2_1__10,
                          linha2_1__9,linha2_1__8,linha2_1__7,linha2_1__6,
                          linha2_1__5,linha2_1__4,linha2_1__3,linha2_1__2,
                          linha2_1__1,linha2_1__0}), .b ({linha3_1__63,
                          linha3_1__62,linha3_1__61,linha3_1__60,linha3_1__59,
                          linha3_1__58,linha3_1__57,linha3_1__56,linha3_1__55,
                          linha3_1__54,linha3_1__53,linha3_1__52,linha3_1__51,
                          linha3_1__50,linha3_1__49,linha3_1__48,linha3_1__47,
                          linha3_1__46,linha3_1__45,linha3_1__44,linha3_1__43,
                          linha3_1__42,linha3_1__41,linha3_1__40,linha3_1__39,
                          linha3_1__38,linha3_1__37,linha3_1__36,linha3_1__35,
                          linha3_1__34,linha3_1__33,linha3_1__32,linha3_1__31,
                          linha3_1__30,linha3_1__29,linha3_1__28,linha3_1__27,
                          linha3_1__26,linha3_1__25,linha3_1__24,linha3_1__23,
                          linha3_1__22,linha3_1__21,linha3_1__20,linha3_1__19,
                          linha3_1__18,linha3_1__17,linha3_1__16,linha3_1__15,
                          linha3_1__14,linha3_1__13,linha3_1__12,linha3_1__11,
                          linha3_1__10,linha3_1__9,linha3_1__8,linha3_1__7,
                          linha3_1__6,linha3_1__5,linha3_1__4,linha3_1__3,
                          linha3_1__2,linha3_1__1,linha3_1__0})) ;
    Mux2x1_64 row_1_rowi_bni1_muxMax (.r ({linha2_2__63,linha2_2__62,
              linha2_2__61,linha2_2__60,linha2_2__59,linha2_2__58,linha2_2__57,
              linha2_2__56,linha2_2__55,linha2_2__54,linha2_2__53,linha2_2__52,
              linha2_2__51,linha2_2__50,linha2_2__49,linha2_2__48,linha2_2__47,
              linha2_2__46,linha2_2__45,linha2_2__44,linha2_2__43,linha2_2__42,
              linha2_2__41,linha2_2__40,linha2_2__39,linha2_2__38,linha2_2__37,
              linha2_2__36,linha2_2__35,linha2_2__34,linha2_2__33,linha2_2__32,
              linha2_2__31,linha2_2__30,linha2_2__29,linha2_2__28,linha2_2__27,
              linha2_2__26,linha2_2__25,linha2_2__24,linha2_2__23,linha2_2__22,
              linha2_2__21,linha2_2__20,linha2_2__19,linha2_2__18,linha2_2__17,
              linha2_2__16,linha2_2__15,linha2_2__14,linha2_2__13,linha2_2__12,
              linha2_2__11,linha2_2__10,linha2_2__9,linha2_2__8,linha2_2__7,
              linha2_2__6,linha2_2__5,linha2_2__4,linha2_2__3,linha2_2__2,
              linha2_2__1,linha2_2__0}), .a1 ({linha3_1__63,linha3_1__62,
              linha3_1__61,linha3_1__60,linha3_1__59,linha3_1__58,linha3_1__57,
              linha3_1__56,linha3_1__55,linha3_1__54,linha3_1__53,linha3_1__52,
              linha3_1__51,linha3_1__50,linha3_1__49,linha3_1__48,linha3_1__47,
              linha3_1__46,linha3_1__45,linha3_1__44,linha3_1__43,linha3_1__42,
              linha3_1__41,linha3_1__40,linha3_1__39,linha3_1__38,linha3_1__37,
              linha3_1__36,linha3_1__35,linha3_1__34,linha3_1__33,linha3_1__32,
              linha3_1__31,linha3_1__30,linha3_1__29,linha3_1__28,linha3_1__27,
              linha3_1__26,linha3_1__25,linha3_1__24,linha3_1__23,linha3_1__22,
              linha3_1__21,linha3_1__20,linha3_1__19,linha3_1__18,linha3_1__17,
              linha3_1__16,linha3_1__15,linha3_1__14,linha3_1__13,linha3_1__12,
              linha3_1__11,linha3_1__10,linha3_1__9,linha3_1__8,linha3_1__7,
              linha3_1__6,linha3_1__5,linha3_1__4,linha3_1__3,linha3_1__2,
              linha3_1__1,linha3_1__0}), .a0 ({linha2_1__63,linha2_1__62,
              linha2_1__61,linha2_1__60,linha2_1__59,linha2_1__58,linha2_1__57,
              linha2_1__56,linha2_1__55,linha2_1__54,linha2_1__53,linha2_1__52,
              linha2_1__51,linha2_1__50,linha2_1__49,linha2_1__48,linha2_1__47,
              linha2_1__46,linha2_1__45,linha2_1__44,linha2_1__43,linha2_1__42,
              linha2_1__41,linha2_1__40,linha2_1__39,linha2_1__38,linha2_1__37,
              linha2_1__36,linha2_1__35,linha2_1__34,linha2_1__33,linha2_1__32,
              linha2_1__31,linha2_1__30,linha2_1__29,linha2_1__28,linha2_1__27,
              linha2_1__26,linha2_1__25,linha2_1__24,linha2_1__23,linha2_1__22,
              linha2_1__21,linha2_1__20,linha2_1__19,linha2_1__18,linha2_1__17,
              linha2_1__16,linha2_1__15,linha2_1__14,linha2_1__13,linha2_1__12,
              linha2_1__11,linha2_1__10,linha2_1__9,linha2_1__8,linha2_1__7,
              linha2_1__6,linha2_1__5,linha2_1__4,linha2_1__3,linha2_1__2,
              linha2_1__1,linha2_1__0}), .s (row_1_rowi_bni1_l)) ;
    Mux2x1_64 row_1_rowi_bni1_muxMin (.r ({linha3_2__63,linha3_2__62,
              linha3_2__61,linha3_2__60,linha3_2__59,linha3_2__58,linha3_2__57,
              linha3_2__56,linha3_2__55,linha3_2__54,linha3_2__53,linha3_2__52,
              linha3_2__51,linha3_2__50,linha3_2__49,linha3_2__48,linha3_2__47,
              linha3_2__46,linha3_2__45,linha3_2__44,linha3_2__43,linha3_2__42,
              linha3_2__41,linha3_2__40,linha3_2__39,linha3_2__38,linha3_2__37,
              linha3_2__36,linha3_2__35,linha3_2__34,linha3_2__33,linha3_2__32,
              linha3_2__31,linha3_2__30,linha3_2__29,linha3_2__28,linha3_2__27,
              linha3_2__26,linha3_2__25,linha3_2__24,linha3_2__23,linha3_2__22,
              linha3_2__21,linha3_2__20,linha3_2__19,linha3_2__18,linha3_2__17,
              linha3_2__16,linha3_2__15,linha3_2__14,linha3_2__13,linha3_2__12,
              linha3_2__11,linha3_2__10,linha3_2__9,linha3_2__8,linha3_2__7,
              linha3_2__6,linha3_2__5,linha3_2__4,linha3_2__3,linha3_2__2,
              linha3_2__1,linha3_2__0}), .a1 ({linha2_1__63,linha2_1__62,
              linha2_1__61,linha2_1__60,linha2_1__59,linha2_1__58,linha2_1__57,
              linha2_1__56,linha2_1__55,linha2_1__54,linha2_1__53,linha2_1__52,
              linha2_1__51,linha2_1__50,linha2_1__49,linha2_1__48,linha2_1__47,
              linha2_1__46,linha2_1__45,linha2_1__44,linha2_1__43,linha2_1__42,
              linha2_1__41,linha2_1__40,linha2_1__39,linha2_1__38,linha2_1__37,
              linha2_1__36,linha2_1__35,linha2_1__34,linha2_1__33,linha2_1__32,
              linha2_1__31,linha2_1__30,linha2_1__29,linha2_1__28,linha2_1__27,
              linha2_1__26,linha2_1__25,linha2_1__24,linha2_1__23,linha2_1__22,
              linha2_1__21,linha2_1__20,linha2_1__19,linha2_1__18,linha2_1__17,
              linha2_1__16,linha2_1__15,linha2_1__14,linha2_1__13,linha2_1__12,
              linha2_1__11,linha2_1__10,linha2_1__9,linha2_1__8,linha2_1__7,
              linha2_1__6,linha2_1__5,linha2_1__4,linha2_1__3,linha2_1__2,
              linha2_1__1,linha2_1__0}), .a0 ({linha3_1__63,linha3_1__62,
              linha3_1__61,linha3_1__60,linha3_1__59,linha3_1__58,linha3_1__57,
              linha3_1__56,linha3_1__55,linha3_1__54,linha3_1__53,linha3_1__52,
              linha3_1__51,linha3_1__50,linha3_1__49,linha3_1__48,linha3_1__47,
              linha3_1__46,linha3_1__45,linha3_1__44,linha3_1__43,linha3_1__42,
              linha3_1__41,linha3_1__40,linha3_1__39,linha3_1__38,linha3_1__37,
              linha3_1__36,linha3_1__35,linha3_1__34,linha3_1__33,linha3_1__32,
              linha3_1__31,linha3_1__30,linha3_1__29,linha3_1__28,linha3_1__27,
              linha3_1__26,linha3_1__25,linha3_1__24,linha3_1__23,linha3_1__22,
              linha3_1__21,linha3_1__20,linha3_1__19,linha3_1__18,linha3_1__17,
              linha3_1__16,linha3_1__15,linha3_1__14,linha3_1__13,linha3_1__12,
              linha3_1__11,linha3_1__10,linha3_1__9,linha3_1__8,linha3_1__7,
              linha3_1__6,linha3_1__5,linha3_1__4,linha3_1__3,linha3_1__2,
              linha3_1__1,linha3_1__0}), .s (row_1_rowi_bni1_l)) ;
    juntarComparadores_64 row_1_rowi_bni2_Comp (.g (\$dummy [5]), .l (
                          row_1_rowi_bni2_l), .a ({linha4_1__63,linha4_1__62,
                          linha4_1__61,linha4_1__60,linha4_1__59,linha4_1__58,
                          linha4_1__57,linha4_1__56,linha4_1__55,linha4_1__54,
                          linha4_1__53,linha4_1__52,linha4_1__51,linha4_1__50,
                          linha4_1__49,linha4_1__48,linha4_1__47,linha4_1__46,
                          linha4_1__45,linha4_1__44,linha4_1__43,linha4_1__42,
                          linha4_1__41,linha4_1__40,linha4_1__39,linha4_1__38,
                          linha4_1__37,linha4_1__36,linha4_1__35,linha4_1__34,
                          linha4_1__33,linha4_1__32,linha4_1__31,linha4_1__30,
                          linha4_1__29,linha4_1__28,linha4_1__27,linha4_1__26,
                          linha4_1__25,linha4_1__24,linha4_1__23,linha4_1__22,
                          linha4_1__21,linha4_1__20,linha4_1__19,linha4_1__18,
                          linha4_1__17,linha4_1__16,linha4_1__15,linha4_1__14,
                          linha4_1__13,linha4_1__12,linha4_1__11,linha4_1__10,
                          linha4_1__9,linha4_1__8,linha4_1__7,linha4_1__6,
                          linha4_1__5,linha4_1__4,linha4_1__3,linha4_1__2,
                          linha4_1__1,linha4_1__0}), .b ({linha5_1__63,
                          linha5_1__62,linha5_1__61,linha5_1__60,linha5_1__59,
                          linha5_1__58,linha5_1__57,linha5_1__56,linha5_1__55,
                          linha5_1__54,linha5_1__53,linha5_1__52,linha5_1__51,
                          linha5_1__50,linha5_1__49,linha5_1__48,linha5_1__47,
                          linha5_1__46,linha5_1__45,linha5_1__44,linha5_1__43,
                          linha5_1__42,linha5_1__41,linha5_1__40,linha5_1__39,
                          linha5_1__38,linha5_1__37,linha5_1__36,linha5_1__35,
                          linha5_1__34,linha5_1__33,linha5_1__32,linha5_1__31,
                          linha5_1__30,linha5_1__29,linha5_1__28,linha5_1__27,
                          linha5_1__26,linha5_1__25,linha5_1__24,linha5_1__23,
                          linha5_1__22,linha5_1__21,linha5_1__20,linha5_1__19,
                          linha5_1__18,linha5_1__17,linha5_1__16,linha5_1__15,
                          linha5_1__14,linha5_1__13,linha5_1__12,linha5_1__11,
                          linha5_1__10,linha5_1__9,linha5_1__8,linha5_1__7,
                          linha5_1__6,linha5_1__5,linha5_1__4,linha5_1__3,
                          linha5_1__2,linha5_1__1,linha5_1__0})) ;
    Mux2x1_64 row_1_rowi_bni2_muxMax (.r ({linha4_2__63,linha4_2__62,
              linha4_2__61,linha4_2__60,linha4_2__59,linha4_2__58,linha4_2__57,
              linha4_2__56,linha4_2__55,linha4_2__54,linha4_2__53,linha4_2__52,
              linha4_2__51,linha4_2__50,linha4_2__49,linha4_2__48,linha4_2__47,
              linha4_2__46,linha4_2__45,linha4_2__44,linha4_2__43,linha4_2__42,
              linha4_2__41,linha4_2__40,linha4_2__39,linha4_2__38,linha4_2__37,
              linha4_2__36,linha4_2__35,linha4_2__34,linha4_2__33,linha4_2__32,
              linha4_2__31,linha4_2__30,linha4_2__29,linha4_2__28,linha4_2__27,
              linha4_2__26,linha4_2__25,linha4_2__24,linha4_2__23,linha4_2__22,
              linha4_2__21,linha4_2__20,linha4_2__19,linha4_2__18,linha4_2__17,
              linha4_2__16,linha4_2__15,linha4_2__14,linha4_2__13,linha4_2__12,
              linha4_2__11,linha4_2__10,linha4_2__9,linha4_2__8,linha4_2__7,
              linha4_2__6,linha4_2__5,linha4_2__4,linha4_2__3,linha4_2__2,
              linha4_2__1,linha4_2__0}), .a1 ({linha5_1__63,linha5_1__62,
              linha5_1__61,linha5_1__60,linha5_1__59,linha5_1__58,linha5_1__57,
              linha5_1__56,linha5_1__55,linha5_1__54,linha5_1__53,linha5_1__52,
              linha5_1__51,linha5_1__50,linha5_1__49,linha5_1__48,linha5_1__47,
              linha5_1__46,linha5_1__45,linha5_1__44,linha5_1__43,linha5_1__42,
              linha5_1__41,linha5_1__40,linha5_1__39,linha5_1__38,linha5_1__37,
              linha5_1__36,linha5_1__35,linha5_1__34,linha5_1__33,linha5_1__32,
              linha5_1__31,linha5_1__30,linha5_1__29,linha5_1__28,linha5_1__27,
              linha5_1__26,linha5_1__25,linha5_1__24,linha5_1__23,linha5_1__22,
              linha5_1__21,linha5_1__20,linha5_1__19,linha5_1__18,linha5_1__17,
              linha5_1__16,linha5_1__15,linha5_1__14,linha5_1__13,linha5_1__12,
              linha5_1__11,linha5_1__10,linha5_1__9,linha5_1__8,linha5_1__7,
              linha5_1__6,linha5_1__5,linha5_1__4,linha5_1__3,linha5_1__2,
              linha5_1__1,linha5_1__0}), .a0 ({linha4_1__63,linha4_1__62,
              linha4_1__61,linha4_1__60,linha4_1__59,linha4_1__58,linha4_1__57,
              linha4_1__56,linha4_1__55,linha4_1__54,linha4_1__53,linha4_1__52,
              linha4_1__51,linha4_1__50,linha4_1__49,linha4_1__48,linha4_1__47,
              linha4_1__46,linha4_1__45,linha4_1__44,linha4_1__43,linha4_1__42,
              linha4_1__41,linha4_1__40,linha4_1__39,linha4_1__38,linha4_1__37,
              linha4_1__36,linha4_1__35,linha4_1__34,linha4_1__33,linha4_1__32,
              linha4_1__31,linha4_1__30,linha4_1__29,linha4_1__28,linha4_1__27,
              linha4_1__26,linha4_1__25,linha4_1__24,linha4_1__23,linha4_1__22,
              linha4_1__21,linha4_1__20,linha4_1__19,linha4_1__18,linha4_1__17,
              linha4_1__16,linha4_1__15,linha4_1__14,linha4_1__13,linha4_1__12,
              linha4_1__11,linha4_1__10,linha4_1__9,linha4_1__8,linha4_1__7,
              linha4_1__6,linha4_1__5,linha4_1__4,linha4_1__3,linha4_1__2,
              linha4_1__1,linha4_1__0}), .s (row_1_rowi_bni2_l)) ;
    Mux2x1_64 row_1_rowi_bni2_muxMin (.r ({linha5_2__63,linha5_2__62,
              linha5_2__61,linha5_2__60,linha5_2__59,linha5_2__58,linha5_2__57,
              linha5_2__56,linha5_2__55,linha5_2__54,linha5_2__53,linha5_2__52,
              linha5_2__51,linha5_2__50,linha5_2__49,linha5_2__48,linha5_2__47,
              linha5_2__46,linha5_2__45,linha5_2__44,linha5_2__43,linha5_2__42,
              linha5_2__41,linha5_2__40,linha5_2__39,linha5_2__38,linha5_2__37,
              linha5_2__36,linha5_2__35,linha5_2__34,linha5_2__33,linha5_2__32,
              linha5_2__31,linha5_2__30,linha5_2__29,linha5_2__28,linha5_2__27,
              linha5_2__26,linha5_2__25,linha5_2__24,linha5_2__23,linha5_2__22,
              linha5_2__21,linha5_2__20,linha5_2__19,linha5_2__18,linha5_2__17,
              linha5_2__16,linha5_2__15,linha5_2__14,linha5_2__13,linha5_2__12,
              linha5_2__11,linha5_2__10,linha5_2__9,linha5_2__8,linha5_2__7,
              linha5_2__6,linha5_2__5,linha5_2__4,linha5_2__3,linha5_2__2,
              linha5_2__1,linha5_2__0}), .a1 ({linha4_1__63,linha4_1__62,
              linha4_1__61,linha4_1__60,linha4_1__59,linha4_1__58,linha4_1__57,
              linha4_1__56,linha4_1__55,linha4_1__54,linha4_1__53,linha4_1__52,
              linha4_1__51,linha4_1__50,linha4_1__49,linha4_1__48,linha4_1__47,
              linha4_1__46,linha4_1__45,linha4_1__44,linha4_1__43,linha4_1__42,
              linha4_1__41,linha4_1__40,linha4_1__39,linha4_1__38,linha4_1__37,
              linha4_1__36,linha4_1__35,linha4_1__34,linha4_1__33,linha4_1__32,
              linha4_1__31,linha4_1__30,linha4_1__29,linha4_1__28,linha4_1__27,
              linha4_1__26,linha4_1__25,linha4_1__24,linha4_1__23,linha4_1__22,
              linha4_1__21,linha4_1__20,linha4_1__19,linha4_1__18,linha4_1__17,
              linha4_1__16,linha4_1__15,linha4_1__14,linha4_1__13,linha4_1__12,
              linha4_1__11,linha4_1__10,linha4_1__9,linha4_1__8,linha4_1__7,
              linha4_1__6,linha4_1__5,linha4_1__4,linha4_1__3,linha4_1__2,
              linha4_1__1,linha4_1__0}), .a0 ({linha5_1__63,linha5_1__62,
              linha5_1__61,linha5_1__60,linha5_1__59,linha5_1__58,linha5_1__57,
              linha5_1__56,linha5_1__55,linha5_1__54,linha5_1__53,linha5_1__52,
              linha5_1__51,linha5_1__50,linha5_1__49,linha5_1__48,linha5_1__47,
              linha5_1__46,linha5_1__45,linha5_1__44,linha5_1__43,linha5_1__42,
              linha5_1__41,linha5_1__40,linha5_1__39,linha5_1__38,linha5_1__37,
              linha5_1__36,linha5_1__35,linha5_1__34,linha5_1__33,linha5_1__32,
              linha5_1__31,linha5_1__30,linha5_1__29,linha5_1__28,linha5_1__27,
              linha5_1__26,linha5_1__25,linha5_1__24,linha5_1__23,linha5_1__22,
              linha5_1__21,linha5_1__20,linha5_1__19,linha5_1__18,linha5_1__17,
              linha5_1__16,linha5_1__15,linha5_1__14,linha5_1__13,linha5_1__12,
              linha5_1__11,linha5_1__10,linha5_1__9,linha5_1__8,linha5_1__7,
              linha5_1__6,linha5_1__5,linha5_1__4,linha5_1__3,linha5_1__2,
              linha5_1__1,linha5_1__0}), .s (row_1_rowi_bni2_l)) ;
    juntarComparadores_64 row_1_rowi_bni3_Comp (.g (\$dummy [6]), .l (
                          row_1_rowi_bni3_l), .a ({linha6_1__63,linha6_1__62,
                          linha6_1__61,linha6_1__60,linha6_1__59,linha6_1__58,
                          linha6_1__57,linha6_1__56,linha6_1__55,linha6_1__54,
                          linha6_1__53,linha6_1__52,linha6_1__51,linha6_1__50,
                          linha6_1__49,linha6_1__48,linha6_1__47,linha6_1__46,
                          linha6_1__45,linha6_1__44,linha6_1__43,linha6_1__42,
                          linha6_1__41,linha6_1__40,linha6_1__39,linha6_1__38,
                          linha6_1__37,linha6_1__36,linha6_1__35,linha6_1__34,
                          linha6_1__33,linha6_1__32,linha6_1__31,linha6_1__30,
                          linha6_1__29,linha6_1__28,linha6_1__27,linha6_1__26,
                          linha6_1__25,linha6_1__24,linha6_1__23,linha6_1__22,
                          linha6_1__21,linha6_1__20,linha6_1__19,linha6_1__18,
                          linha6_1__17,linha6_1__16,linha6_1__15,linha6_1__14,
                          linha6_1__13,linha6_1__12,linha6_1__11,linha6_1__10,
                          linha6_1__9,linha6_1__8,linha6_1__7,linha6_1__6,
                          linha6_1__5,linha6_1__4,linha6_1__3,linha6_1__2,
                          linha6_1__1,linha6_1__0}), .b ({linha7_1__63,
                          linha7_1__62,linha7_1__61,linha7_1__60,linha7_1__59,
                          linha7_1__58,linha7_1__57,linha7_1__56,linha7_1__55,
                          linha7_1__54,linha7_1__53,linha7_1__52,linha7_1__51,
                          linha7_1__50,linha7_1__49,linha7_1__48,linha7_1__47,
                          linha7_1__46,linha7_1__45,linha7_1__44,linha7_1__43,
                          linha7_1__42,linha7_1__41,linha7_1__40,linha7_1__39,
                          linha7_1__38,linha7_1__37,linha7_1__36,linha7_1__35,
                          linha7_1__34,linha7_1__33,linha7_1__32,linha7_1__31,
                          linha7_1__30,linha7_1__29,linha7_1__28,linha7_1__27,
                          linha7_1__26,linha7_1__25,linha7_1__24,linha7_1__23,
                          linha7_1__22,linha7_1__21,linha7_1__20,linha7_1__19,
                          linha7_1__18,linha7_1__17,linha7_1__16,linha7_1__15,
                          linha7_1__14,linha7_1__13,linha7_1__12,linha7_1__11,
                          linha7_1__10,linha7_1__9,linha7_1__8,linha7_1__7,
                          linha7_1__6,linha7_1__5,linha7_1__4,linha7_1__3,
                          linha7_1__2,linha7_1__1,linha7_1__0})) ;
    Mux2x1_64 row_1_rowi_bni3_muxMax (.r ({linha6_2__63,linha6_2__62,
              linha6_2__61,linha6_2__60,linha6_2__59,linha6_2__58,linha6_2__57,
              linha6_2__56,linha6_2__55,linha6_2__54,linha6_2__53,linha6_2__52,
              linha6_2__51,linha6_2__50,linha6_2__49,linha6_2__48,linha6_2__47,
              linha6_2__46,linha6_2__45,linha6_2__44,linha6_2__43,linha6_2__42,
              linha6_2__41,linha6_2__40,linha6_2__39,linha6_2__38,linha6_2__37,
              linha6_2__36,linha6_2__35,linha6_2__34,linha6_2__33,linha6_2__32,
              linha6_2__31,linha6_2__30,linha6_2__29,linha6_2__28,linha6_2__27,
              linha6_2__26,linha6_2__25,linha6_2__24,linha6_2__23,linha6_2__22,
              linha6_2__21,linha6_2__20,linha6_2__19,linha6_2__18,linha6_2__17,
              linha6_2__16,linha6_2__15,linha6_2__14,linha6_2__13,linha6_2__12,
              linha6_2__11,linha6_2__10,linha6_2__9,linha6_2__8,linha6_2__7,
              linha6_2__6,linha6_2__5,linha6_2__4,linha6_2__3,linha6_2__2,
              linha6_2__1,linha6_2__0}), .a1 ({linha7_1__63,linha7_1__62,
              linha7_1__61,linha7_1__60,linha7_1__59,linha7_1__58,linha7_1__57,
              linha7_1__56,linha7_1__55,linha7_1__54,linha7_1__53,linha7_1__52,
              linha7_1__51,linha7_1__50,linha7_1__49,linha7_1__48,linha7_1__47,
              linha7_1__46,linha7_1__45,linha7_1__44,linha7_1__43,linha7_1__42,
              linha7_1__41,linha7_1__40,linha7_1__39,linha7_1__38,linha7_1__37,
              linha7_1__36,linha7_1__35,linha7_1__34,linha7_1__33,linha7_1__32,
              linha7_1__31,linha7_1__30,linha7_1__29,linha7_1__28,linha7_1__27,
              linha7_1__26,linha7_1__25,linha7_1__24,linha7_1__23,linha7_1__22,
              linha7_1__21,linha7_1__20,linha7_1__19,linha7_1__18,linha7_1__17,
              linha7_1__16,linha7_1__15,linha7_1__14,linha7_1__13,linha7_1__12,
              linha7_1__11,linha7_1__10,linha7_1__9,linha7_1__8,linha7_1__7,
              linha7_1__6,linha7_1__5,linha7_1__4,linha7_1__3,linha7_1__2,
              linha7_1__1,linha7_1__0}), .a0 ({linha6_1__63,linha6_1__62,
              linha6_1__61,linha6_1__60,linha6_1__59,linha6_1__58,linha6_1__57,
              linha6_1__56,linha6_1__55,linha6_1__54,linha6_1__53,linha6_1__52,
              linha6_1__51,linha6_1__50,linha6_1__49,linha6_1__48,linha6_1__47,
              linha6_1__46,linha6_1__45,linha6_1__44,linha6_1__43,linha6_1__42,
              linha6_1__41,linha6_1__40,linha6_1__39,linha6_1__38,linha6_1__37,
              linha6_1__36,linha6_1__35,linha6_1__34,linha6_1__33,linha6_1__32,
              linha6_1__31,linha6_1__30,linha6_1__29,linha6_1__28,linha6_1__27,
              linha6_1__26,linha6_1__25,linha6_1__24,linha6_1__23,linha6_1__22,
              linha6_1__21,linha6_1__20,linha6_1__19,linha6_1__18,linha6_1__17,
              linha6_1__16,linha6_1__15,linha6_1__14,linha6_1__13,linha6_1__12,
              linha6_1__11,linha6_1__10,linha6_1__9,linha6_1__8,linha6_1__7,
              linha6_1__6,linha6_1__5,linha6_1__4,linha6_1__3,linha6_1__2,
              linha6_1__1,linha6_1__0}), .s (row_1_rowi_bni3_l)) ;
    Mux2x1_64 row_1_rowi_bni3_muxMin (.r ({linha7_2__63,linha7_2__62,
              linha7_2__61,linha7_2__60,linha7_2__59,linha7_2__58,linha7_2__57,
              linha7_2__56,linha7_2__55,linha7_2__54,linha7_2__53,linha7_2__52,
              linha7_2__51,linha7_2__50,linha7_2__49,linha7_2__48,linha7_2__47,
              linha7_2__46,linha7_2__45,linha7_2__44,linha7_2__43,linha7_2__42,
              linha7_2__41,linha7_2__40,linha7_2__39,linha7_2__38,linha7_2__37,
              linha7_2__36,linha7_2__35,linha7_2__34,linha7_2__33,linha7_2__32,
              linha7_2__31,linha7_2__30,linha7_2__29,linha7_2__28,linha7_2__27,
              linha7_2__26,linha7_2__25,linha7_2__24,linha7_2__23,linha7_2__22,
              linha7_2__21,linha7_2__20,linha7_2__19,linha7_2__18,linha7_2__17,
              linha7_2__16,linha7_2__15,linha7_2__14,linha7_2__13,linha7_2__12,
              linha7_2__11,linha7_2__10,linha7_2__9,linha7_2__8,linha7_2__7,
              linha7_2__6,linha7_2__5,linha7_2__4,linha7_2__3,linha7_2__2,
              linha7_2__1,linha7_2__0}), .a1 ({linha6_1__63,linha6_1__62,
              linha6_1__61,linha6_1__60,linha6_1__59,linha6_1__58,linha6_1__57,
              linha6_1__56,linha6_1__55,linha6_1__54,linha6_1__53,linha6_1__52,
              linha6_1__51,linha6_1__50,linha6_1__49,linha6_1__48,linha6_1__47,
              linha6_1__46,linha6_1__45,linha6_1__44,linha6_1__43,linha6_1__42,
              linha6_1__41,linha6_1__40,linha6_1__39,linha6_1__38,linha6_1__37,
              linha6_1__36,linha6_1__35,linha6_1__34,linha6_1__33,linha6_1__32,
              linha6_1__31,linha6_1__30,linha6_1__29,linha6_1__28,linha6_1__27,
              linha6_1__26,linha6_1__25,linha6_1__24,linha6_1__23,linha6_1__22,
              linha6_1__21,linha6_1__20,linha6_1__19,linha6_1__18,linha6_1__17,
              linha6_1__16,linha6_1__15,linha6_1__14,linha6_1__13,linha6_1__12,
              linha6_1__11,linha6_1__10,linha6_1__9,linha6_1__8,linha6_1__7,
              linha6_1__6,linha6_1__5,linha6_1__4,linha6_1__3,linha6_1__2,
              linha6_1__1,linha6_1__0}), .a0 ({linha7_1__63,linha7_1__62,
              linha7_1__61,linha7_1__60,linha7_1__59,linha7_1__58,linha7_1__57,
              linha7_1__56,linha7_1__55,linha7_1__54,linha7_1__53,linha7_1__52,
              linha7_1__51,linha7_1__50,linha7_1__49,linha7_1__48,linha7_1__47,
              linha7_1__46,linha7_1__45,linha7_1__44,linha7_1__43,linha7_1__42,
              linha7_1__41,linha7_1__40,linha7_1__39,linha7_1__38,linha7_1__37,
              linha7_1__36,linha7_1__35,linha7_1__34,linha7_1__33,linha7_1__32,
              linha7_1__31,linha7_1__30,linha7_1__29,linha7_1__28,linha7_1__27,
              linha7_1__26,linha7_1__25,linha7_1__24,linha7_1__23,linha7_1__22,
              linha7_1__21,linha7_1__20,linha7_1__19,linha7_1__18,linha7_1__17,
              linha7_1__16,linha7_1__15,linha7_1__14,linha7_1__13,linha7_1__12,
              linha7_1__11,linha7_1__10,linha7_1__9,linha7_1__8,linha7_1__7,
              linha7_1__6,linha7_1__5,linha7_1__4,linha7_1__3,linha7_1__2,
              linha7_1__1,linha7_1__0}), .s (row_1_rowi_bni3_l)) ;
    juntarComparadores_64 row_2_rowp_bni1_Comp (.g (\$dummy [7]), .l (
                          row_2_rowp_bni1_l), .a ({linha1_1__63,linha1_1__62,
                          linha1_1__61,linha1_1__60,linha1_1__59,linha1_1__58,
                          linha1_1__57,linha1_1__56,linha1_1__55,linha1_1__54,
                          linha1_1__53,linha1_1__52,linha1_1__51,linha1_1__50,
                          linha1_1__49,linha1_1__48,linha1_1__47,linha1_1__46,
                          linha1_1__45,linha1_1__44,linha1_1__43,linha1_1__42,
                          linha1_1__41,linha1_1__40,linha1_1__39,linha1_1__38,
                          linha1_1__37,linha1_1__36,linha1_1__35,linha1_1__34,
                          linha1_1__33,linha1_1__32,linha1_1__31,linha1_1__30,
                          linha1_1__29,linha1_1__28,linha1_1__27,linha1_1__26,
                          linha1_1__25,linha1_1__24,linha1_1__23,linha1_1__22,
                          linha1_1__21,linha1_1__20,linha1_1__19,linha1_1__18,
                          linha1_1__17,linha1_1__16,linha1_1__15,linha1_1__14,
                          linha1_1__13,linha1_1__12,linha1_1__11,linha1_1__10,
                          linha1_1__9,linha1_1__8,linha1_1__7,linha1_1__6,
                          linha1_1__5,linha1_1__4,linha1_1__3,linha1_1__2,
                          linha1_1__1,linha1_1__0}), .b ({linha2_2__63,
                          linha2_2__62,linha2_2__61,linha2_2__60,linha2_2__59,
                          linha2_2__58,linha2_2__57,linha2_2__56,linha2_2__55,
                          linha2_2__54,linha2_2__53,linha2_2__52,linha2_2__51,
                          linha2_2__50,linha2_2__49,linha2_2__48,linha2_2__47,
                          linha2_2__46,linha2_2__45,linha2_2__44,linha2_2__43,
                          linha2_2__42,linha2_2__41,linha2_2__40,linha2_2__39,
                          linha2_2__38,linha2_2__37,linha2_2__36,linha2_2__35,
                          linha2_2__34,linha2_2__33,linha2_2__32,linha2_2__31,
                          linha2_2__30,linha2_2__29,linha2_2__28,linha2_2__27,
                          linha2_2__26,linha2_2__25,linha2_2__24,linha2_2__23,
                          linha2_2__22,linha2_2__21,linha2_2__20,linha2_2__19,
                          linha2_2__18,linha2_2__17,linha2_2__16,linha2_2__15,
                          linha2_2__14,linha2_2__13,linha2_2__12,linha2_2__11,
                          linha2_2__10,linha2_2__9,linha2_2__8,linha2_2__7,
                          linha2_2__6,linha2_2__5,linha2_2__4,linha2_2__3,
                          linha2_2__2,linha2_2__1,linha2_2__0})) ;
    Mux2x1_64 row_2_rowp_bni1_muxMax (.r ({linha1_2__63,linha1_2__62,
              linha1_2__61,linha1_2__60,linha1_2__59,linha1_2__58,linha1_2__57,
              linha1_2__56,linha1_2__55,linha1_2__54,linha1_2__53,linha1_2__52,
              linha1_2__51,linha1_2__50,linha1_2__49,linha1_2__48,linha1_2__47,
              linha1_2__46,linha1_2__45,linha1_2__44,linha1_2__43,linha1_2__42,
              linha1_2__41,linha1_2__40,linha1_2__39,linha1_2__38,linha1_2__37,
              linha1_2__36,linha1_2__35,linha1_2__34,linha1_2__33,linha1_2__32,
              linha1_2__31,linha1_2__30,linha1_2__29,linha1_2__28,linha1_2__27,
              linha1_2__26,linha1_2__25,linha1_2__24,linha1_2__23,linha1_2__22,
              linha1_2__21,linha1_2__20,linha1_2__19,linha1_2__18,linha1_2__17,
              linha1_2__16,linha1_2__15,linha1_2__14,linha1_2__13,linha1_2__12,
              linha1_2__11,linha1_2__10,linha1_2__9,linha1_2__8,linha1_2__7,
              linha1_2__6,linha1_2__5,linha1_2__4,linha1_2__3,linha1_2__2,
              linha1_2__1,linha1_2__0}), .a1 ({linha2_2__63,linha2_2__62,
              linha2_2__61,linha2_2__60,linha2_2__59,linha2_2__58,linha2_2__57,
              linha2_2__56,linha2_2__55,linha2_2__54,linha2_2__53,linha2_2__52,
              linha2_2__51,linha2_2__50,linha2_2__49,linha2_2__48,linha2_2__47,
              linha2_2__46,linha2_2__45,linha2_2__44,linha2_2__43,linha2_2__42,
              linha2_2__41,linha2_2__40,linha2_2__39,linha2_2__38,linha2_2__37,
              linha2_2__36,linha2_2__35,linha2_2__34,linha2_2__33,linha2_2__32,
              linha2_2__31,linha2_2__30,linha2_2__29,linha2_2__28,linha2_2__27,
              linha2_2__26,linha2_2__25,linha2_2__24,linha2_2__23,linha2_2__22,
              linha2_2__21,linha2_2__20,linha2_2__19,linha2_2__18,linha2_2__17,
              linha2_2__16,linha2_2__15,linha2_2__14,linha2_2__13,linha2_2__12,
              linha2_2__11,linha2_2__10,linha2_2__9,linha2_2__8,linha2_2__7,
              linha2_2__6,linha2_2__5,linha2_2__4,linha2_2__3,linha2_2__2,
              linha2_2__1,linha2_2__0}), .a0 ({linha1_1__63,linha1_1__62,
              linha1_1__61,linha1_1__60,linha1_1__59,linha1_1__58,linha1_1__57,
              linha1_1__56,linha1_1__55,linha1_1__54,linha1_1__53,linha1_1__52,
              linha1_1__51,linha1_1__50,linha1_1__49,linha1_1__48,linha1_1__47,
              linha1_1__46,linha1_1__45,linha1_1__44,linha1_1__43,linha1_1__42,
              linha1_1__41,linha1_1__40,linha1_1__39,linha1_1__38,linha1_1__37,
              linha1_1__36,linha1_1__35,linha1_1__34,linha1_1__33,linha1_1__32,
              linha1_1__31,linha1_1__30,linha1_1__29,linha1_1__28,linha1_1__27,
              linha1_1__26,linha1_1__25,linha1_1__24,linha1_1__23,linha1_1__22,
              linha1_1__21,linha1_1__20,linha1_1__19,linha1_1__18,linha1_1__17,
              linha1_1__16,linha1_1__15,linha1_1__14,linha1_1__13,linha1_1__12,
              linha1_1__11,linha1_1__10,linha1_1__9,linha1_1__8,linha1_1__7,
              linha1_1__6,linha1_1__5,linha1_1__4,linha1_1__3,linha1_1__2,
              linha1_1__1,linha1_1__0}), .s (row_2_rowp_bni1_l)) ;
    Mux2x1_64 row_2_rowp_bni1_muxMin (.r ({linha2_3__63,linha2_3__62,
              linha2_3__61,linha2_3__60,linha2_3__59,linha2_3__58,linha2_3__57,
              linha2_3__56,linha2_3__55,linha2_3__54,linha2_3__53,linha2_3__52,
              linha2_3__51,linha2_3__50,linha2_3__49,linha2_3__48,linha2_3__47,
              linha2_3__46,linha2_3__45,linha2_3__44,linha2_3__43,linha2_3__42,
              linha2_3__41,linha2_3__40,linha2_3__39,linha2_3__38,linha2_3__37,
              linha2_3__36,linha2_3__35,linha2_3__34,linha2_3__33,linha2_3__32,
              linha2_3__31,linha2_3__30,linha2_3__29,linha2_3__28,linha2_3__27,
              linha2_3__26,linha2_3__25,linha2_3__24,linha2_3__23,linha2_3__22,
              linha2_3__21,linha2_3__20,linha2_3__19,linha2_3__18,linha2_3__17,
              linha2_3__16,linha2_3__15,linha2_3__14,linha2_3__13,linha2_3__12,
              linha2_3__11,linha2_3__10,linha2_3__9,linha2_3__8,linha2_3__7,
              linha2_3__6,linha2_3__5,linha2_3__4,linha2_3__3,linha2_3__2,
              linha2_3__1,linha2_3__0}), .a1 ({linha1_1__63,linha1_1__62,
              linha1_1__61,linha1_1__60,linha1_1__59,linha1_1__58,linha1_1__57,
              linha1_1__56,linha1_1__55,linha1_1__54,linha1_1__53,linha1_1__52,
              linha1_1__51,linha1_1__50,linha1_1__49,linha1_1__48,linha1_1__47,
              linha1_1__46,linha1_1__45,linha1_1__44,linha1_1__43,linha1_1__42,
              linha1_1__41,linha1_1__40,linha1_1__39,linha1_1__38,linha1_1__37,
              linha1_1__36,linha1_1__35,linha1_1__34,linha1_1__33,linha1_1__32,
              linha1_1__31,linha1_1__30,linha1_1__29,linha1_1__28,linha1_1__27,
              linha1_1__26,linha1_1__25,linha1_1__24,linha1_1__23,linha1_1__22,
              linha1_1__21,linha1_1__20,linha1_1__19,linha1_1__18,linha1_1__17,
              linha1_1__16,linha1_1__15,linha1_1__14,linha1_1__13,linha1_1__12,
              linha1_1__11,linha1_1__10,linha1_1__9,linha1_1__8,linha1_1__7,
              linha1_1__6,linha1_1__5,linha1_1__4,linha1_1__3,linha1_1__2,
              linha1_1__1,linha1_1__0}), .a0 ({linha2_2__63,linha2_2__62,
              linha2_2__61,linha2_2__60,linha2_2__59,linha2_2__58,linha2_2__57,
              linha2_2__56,linha2_2__55,linha2_2__54,linha2_2__53,linha2_2__52,
              linha2_2__51,linha2_2__50,linha2_2__49,linha2_2__48,linha2_2__47,
              linha2_2__46,linha2_2__45,linha2_2__44,linha2_2__43,linha2_2__42,
              linha2_2__41,linha2_2__40,linha2_2__39,linha2_2__38,linha2_2__37,
              linha2_2__36,linha2_2__35,linha2_2__34,linha2_2__33,linha2_2__32,
              linha2_2__31,linha2_2__30,linha2_2__29,linha2_2__28,linha2_2__27,
              linha2_2__26,linha2_2__25,linha2_2__24,linha2_2__23,linha2_2__22,
              linha2_2__21,linha2_2__20,linha2_2__19,linha2_2__18,linha2_2__17,
              linha2_2__16,linha2_2__15,linha2_2__14,linha2_2__13,linha2_2__12,
              linha2_2__11,linha2_2__10,linha2_2__9,linha2_2__8,linha2_2__7,
              linha2_2__6,linha2_2__5,linha2_2__4,linha2_2__3,linha2_2__2,
              linha2_2__1,linha2_2__0}), .s (row_2_rowp_bni1_l)) ;
    juntarComparadores_64 row_2_rowp_bni2_Comp (.g (\$dummy [8]), .l (
                          row_2_rowp_bni2_l), .a ({linha3_2__63,linha3_2__62,
                          linha3_2__61,linha3_2__60,linha3_2__59,linha3_2__58,
                          linha3_2__57,linha3_2__56,linha3_2__55,linha3_2__54,
                          linha3_2__53,linha3_2__52,linha3_2__51,linha3_2__50,
                          linha3_2__49,linha3_2__48,linha3_2__47,linha3_2__46,
                          linha3_2__45,linha3_2__44,linha3_2__43,linha3_2__42,
                          linha3_2__41,linha3_2__40,linha3_2__39,linha3_2__38,
                          linha3_2__37,linha3_2__36,linha3_2__35,linha3_2__34,
                          linha3_2__33,linha3_2__32,linha3_2__31,linha3_2__30,
                          linha3_2__29,linha3_2__28,linha3_2__27,linha3_2__26,
                          linha3_2__25,linha3_2__24,linha3_2__23,linha3_2__22,
                          linha3_2__21,linha3_2__20,linha3_2__19,linha3_2__18,
                          linha3_2__17,linha3_2__16,linha3_2__15,linha3_2__14,
                          linha3_2__13,linha3_2__12,linha3_2__11,linha3_2__10,
                          linha3_2__9,linha3_2__8,linha3_2__7,linha3_2__6,
                          linha3_2__5,linha3_2__4,linha3_2__3,linha3_2__2,
                          linha3_2__1,linha3_2__0}), .b ({linha4_2__63,
                          linha4_2__62,linha4_2__61,linha4_2__60,linha4_2__59,
                          linha4_2__58,linha4_2__57,linha4_2__56,linha4_2__55,
                          linha4_2__54,linha4_2__53,linha4_2__52,linha4_2__51,
                          linha4_2__50,linha4_2__49,linha4_2__48,linha4_2__47,
                          linha4_2__46,linha4_2__45,linha4_2__44,linha4_2__43,
                          linha4_2__42,linha4_2__41,linha4_2__40,linha4_2__39,
                          linha4_2__38,linha4_2__37,linha4_2__36,linha4_2__35,
                          linha4_2__34,linha4_2__33,linha4_2__32,linha4_2__31,
                          linha4_2__30,linha4_2__29,linha4_2__28,linha4_2__27,
                          linha4_2__26,linha4_2__25,linha4_2__24,linha4_2__23,
                          linha4_2__22,linha4_2__21,linha4_2__20,linha4_2__19,
                          linha4_2__18,linha4_2__17,linha4_2__16,linha4_2__15,
                          linha4_2__14,linha4_2__13,linha4_2__12,linha4_2__11,
                          linha4_2__10,linha4_2__9,linha4_2__8,linha4_2__7,
                          linha4_2__6,linha4_2__5,linha4_2__4,linha4_2__3,
                          linha4_2__2,linha4_2__1,linha4_2__0})) ;
    Mux2x1_64 row_2_rowp_bni2_muxMax (.r ({linha3_3__63,linha3_3__62,
              linha3_3__61,linha3_3__60,linha3_3__59,linha3_3__58,linha3_3__57,
              linha3_3__56,linha3_3__55,linha3_3__54,linha3_3__53,linha3_3__52,
              linha3_3__51,linha3_3__50,linha3_3__49,linha3_3__48,linha3_3__47,
              linha3_3__46,linha3_3__45,linha3_3__44,linha3_3__43,linha3_3__42,
              linha3_3__41,linha3_3__40,linha3_3__39,linha3_3__38,linha3_3__37,
              linha3_3__36,linha3_3__35,linha3_3__34,linha3_3__33,linha3_3__32,
              linha3_3__31,linha3_3__30,linha3_3__29,linha3_3__28,linha3_3__27,
              linha3_3__26,linha3_3__25,linha3_3__24,linha3_3__23,linha3_3__22,
              linha3_3__21,linha3_3__20,linha3_3__19,linha3_3__18,linha3_3__17,
              linha3_3__16,linha3_3__15,linha3_3__14,linha3_3__13,linha3_3__12,
              linha3_3__11,linha3_3__10,linha3_3__9,linha3_3__8,linha3_3__7,
              linha3_3__6,linha3_3__5,linha3_3__4,linha3_3__3,linha3_3__2,
              linha3_3__1,linha3_3__0}), .a1 ({linha4_2__63,linha4_2__62,
              linha4_2__61,linha4_2__60,linha4_2__59,linha4_2__58,linha4_2__57,
              linha4_2__56,linha4_2__55,linha4_2__54,linha4_2__53,linha4_2__52,
              linha4_2__51,linha4_2__50,linha4_2__49,linha4_2__48,linha4_2__47,
              linha4_2__46,linha4_2__45,linha4_2__44,linha4_2__43,linha4_2__42,
              linha4_2__41,linha4_2__40,linha4_2__39,linha4_2__38,linha4_2__37,
              linha4_2__36,linha4_2__35,linha4_2__34,linha4_2__33,linha4_2__32,
              linha4_2__31,linha4_2__30,linha4_2__29,linha4_2__28,linha4_2__27,
              linha4_2__26,linha4_2__25,linha4_2__24,linha4_2__23,linha4_2__22,
              linha4_2__21,linha4_2__20,linha4_2__19,linha4_2__18,linha4_2__17,
              linha4_2__16,linha4_2__15,linha4_2__14,linha4_2__13,linha4_2__12,
              linha4_2__11,linha4_2__10,linha4_2__9,linha4_2__8,linha4_2__7,
              linha4_2__6,linha4_2__5,linha4_2__4,linha4_2__3,linha4_2__2,
              linha4_2__1,linha4_2__0}), .a0 ({linha3_2__63,linha3_2__62,
              linha3_2__61,linha3_2__60,linha3_2__59,linha3_2__58,linha3_2__57,
              linha3_2__56,linha3_2__55,linha3_2__54,linha3_2__53,linha3_2__52,
              linha3_2__51,linha3_2__50,linha3_2__49,linha3_2__48,linha3_2__47,
              linha3_2__46,linha3_2__45,linha3_2__44,linha3_2__43,linha3_2__42,
              linha3_2__41,linha3_2__40,linha3_2__39,linha3_2__38,linha3_2__37,
              linha3_2__36,linha3_2__35,linha3_2__34,linha3_2__33,linha3_2__32,
              linha3_2__31,linha3_2__30,linha3_2__29,linha3_2__28,linha3_2__27,
              linha3_2__26,linha3_2__25,linha3_2__24,linha3_2__23,linha3_2__22,
              linha3_2__21,linha3_2__20,linha3_2__19,linha3_2__18,linha3_2__17,
              linha3_2__16,linha3_2__15,linha3_2__14,linha3_2__13,linha3_2__12,
              linha3_2__11,linha3_2__10,linha3_2__9,linha3_2__8,linha3_2__7,
              linha3_2__6,linha3_2__5,linha3_2__4,linha3_2__3,linha3_2__2,
              linha3_2__1,linha3_2__0}), .s (row_2_rowp_bni2_l)) ;
    Mux2x1_64 row_2_rowp_bni2_muxMin (.r ({linha4_3__63,linha4_3__62,
              linha4_3__61,linha4_3__60,linha4_3__59,linha4_3__58,linha4_3__57,
              linha4_3__56,linha4_3__55,linha4_3__54,linha4_3__53,linha4_3__52,
              linha4_3__51,linha4_3__50,linha4_3__49,linha4_3__48,linha4_3__47,
              linha4_3__46,linha4_3__45,linha4_3__44,linha4_3__43,linha4_3__42,
              linha4_3__41,linha4_3__40,linha4_3__39,linha4_3__38,linha4_3__37,
              linha4_3__36,linha4_3__35,linha4_3__34,linha4_3__33,linha4_3__32,
              linha4_3__31,linha4_3__30,linha4_3__29,linha4_3__28,linha4_3__27,
              linha4_3__26,linha4_3__25,linha4_3__24,linha4_3__23,linha4_3__22,
              linha4_3__21,linha4_3__20,linha4_3__19,linha4_3__18,linha4_3__17,
              linha4_3__16,linha4_3__15,linha4_3__14,linha4_3__13,linha4_3__12,
              linha4_3__11,linha4_3__10,linha4_3__9,linha4_3__8,linha4_3__7,
              linha4_3__6,linha4_3__5,linha4_3__4,linha4_3__3,linha4_3__2,
              linha4_3__1,linha4_3__0}), .a1 ({linha3_2__63,linha3_2__62,
              linha3_2__61,linha3_2__60,linha3_2__59,linha3_2__58,linha3_2__57,
              linha3_2__56,linha3_2__55,linha3_2__54,linha3_2__53,linha3_2__52,
              linha3_2__51,linha3_2__50,linha3_2__49,linha3_2__48,linha3_2__47,
              linha3_2__46,linha3_2__45,linha3_2__44,linha3_2__43,linha3_2__42,
              linha3_2__41,linha3_2__40,linha3_2__39,linha3_2__38,linha3_2__37,
              linha3_2__36,linha3_2__35,linha3_2__34,linha3_2__33,linha3_2__32,
              linha3_2__31,linha3_2__30,linha3_2__29,linha3_2__28,linha3_2__27,
              linha3_2__26,linha3_2__25,linha3_2__24,linha3_2__23,linha3_2__22,
              linha3_2__21,linha3_2__20,linha3_2__19,linha3_2__18,linha3_2__17,
              linha3_2__16,linha3_2__15,linha3_2__14,linha3_2__13,linha3_2__12,
              linha3_2__11,linha3_2__10,linha3_2__9,linha3_2__8,linha3_2__7,
              linha3_2__6,linha3_2__5,linha3_2__4,linha3_2__3,linha3_2__2,
              linha3_2__1,linha3_2__0}), .a0 ({linha4_2__63,linha4_2__62,
              linha4_2__61,linha4_2__60,linha4_2__59,linha4_2__58,linha4_2__57,
              linha4_2__56,linha4_2__55,linha4_2__54,linha4_2__53,linha4_2__52,
              linha4_2__51,linha4_2__50,linha4_2__49,linha4_2__48,linha4_2__47,
              linha4_2__46,linha4_2__45,linha4_2__44,linha4_2__43,linha4_2__42,
              linha4_2__41,linha4_2__40,linha4_2__39,linha4_2__38,linha4_2__37,
              linha4_2__36,linha4_2__35,linha4_2__34,linha4_2__33,linha4_2__32,
              linha4_2__31,linha4_2__30,linha4_2__29,linha4_2__28,linha4_2__27,
              linha4_2__26,linha4_2__25,linha4_2__24,linha4_2__23,linha4_2__22,
              linha4_2__21,linha4_2__20,linha4_2__19,linha4_2__18,linha4_2__17,
              linha4_2__16,linha4_2__15,linha4_2__14,linha4_2__13,linha4_2__12,
              linha4_2__11,linha4_2__10,linha4_2__9,linha4_2__8,linha4_2__7,
              linha4_2__6,linha4_2__5,linha4_2__4,linha4_2__3,linha4_2__2,
              linha4_2__1,linha4_2__0}), .s (row_2_rowp_bni2_l)) ;
    juntarComparadores_64 row_2_rowp_bni3_Comp (.g (\$dummy [9]), .l (
                          row_2_rowp_bni3_l), .a ({linha5_2__63,linha5_2__62,
                          linha5_2__61,linha5_2__60,linha5_2__59,linha5_2__58,
                          linha5_2__57,linha5_2__56,linha5_2__55,linha5_2__54,
                          linha5_2__53,linha5_2__52,linha5_2__51,linha5_2__50,
                          linha5_2__49,linha5_2__48,linha5_2__47,linha5_2__46,
                          linha5_2__45,linha5_2__44,linha5_2__43,linha5_2__42,
                          linha5_2__41,linha5_2__40,linha5_2__39,linha5_2__38,
                          linha5_2__37,linha5_2__36,linha5_2__35,linha5_2__34,
                          linha5_2__33,linha5_2__32,linha5_2__31,linha5_2__30,
                          linha5_2__29,linha5_2__28,linha5_2__27,linha5_2__26,
                          linha5_2__25,linha5_2__24,linha5_2__23,linha5_2__22,
                          linha5_2__21,linha5_2__20,linha5_2__19,linha5_2__18,
                          linha5_2__17,linha5_2__16,linha5_2__15,linha5_2__14,
                          linha5_2__13,linha5_2__12,linha5_2__11,linha5_2__10,
                          linha5_2__9,linha5_2__8,linha5_2__7,linha5_2__6,
                          linha5_2__5,linha5_2__4,linha5_2__3,linha5_2__2,
                          linha5_2__1,linha5_2__0}), .b ({linha6_2__63,
                          linha6_2__62,linha6_2__61,linha6_2__60,linha6_2__59,
                          linha6_2__58,linha6_2__57,linha6_2__56,linha6_2__55,
                          linha6_2__54,linha6_2__53,linha6_2__52,linha6_2__51,
                          linha6_2__50,linha6_2__49,linha6_2__48,linha6_2__47,
                          linha6_2__46,linha6_2__45,linha6_2__44,linha6_2__43,
                          linha6_2__42,linha6_2__41,linha6_2__40,linha6_2__39,
                          linha6_2__38,linha6_2__37,linha6_2__36,linha6_2__35,
                          linha6_2__34,linha6_2__33,linha6_2__32,linha6_2__31,
                          linha6_2__30,linha6_2__29,linha6_2__28,linha6_2__27,
                          linha6_2__26,linha6_2__25,linha6_2__24,linha6_2__23,
                          linha6_2__22,linha6_2__21,linha6_2__20,linha6_2__19,
                          linha6_2__18,linha6_2__17,linha6_2__16,linha6_2__15,
                          linha6_2__14,linha6_2__13,linha6_2__12,linha6_2__11,
                          linha6_2__10,linha6_2__9,linha6_2__8,linha6_2__7,
                          linha6_2__6,linha6_2__5,linha6_2__4,linha6_2__3,
                          linha6_2__2,linha6_2__1,linha6_2__0})) ;
    Mux2x1_64 row_2_rowp_bni3_muxMax (.r ({linha5_3__63,linha5_3__62,
              linha5_3__61,linha5_3__60,linha5_3__59,linha5_3__58,linha5_3__57,
              linha5_3__56,linha5_3__55,linha5_3__54,linha5_3__53,linha5_3__52,
              linha5_3__51,linha5_3__50,linha5_3__49,linha5_3__48,linha5_3__47,
              linha5_3__46,linha5_3__45,linha5_3__44,linha5_3__43,linha5_3__42,
              linha5_3__41,linha5_3__40,linha5_3__39,linha5_3__38,linha5_3__37,
              linha5_3__36,linha5_3__35,linha5_3__34,linha5_3__33,linha5_3__32,
              linha5_3__31,linha5_3__30,linha5_3__29,linha5_3__28,linha5_3__27,
              linha5_3__26,linha5_3__25,linha5_3__24,linha5_3__23,linha5_3__22,
              linha5_3__21,linha5_3__20,linha5_3__19,linha5_3__18,linha5_3__17,
              linha5_3__16,linha5_3__15,linha5_3__14,linha5_3__13,linha5_3__12,
              linha5_3__11,linha5_3__10,linha5_3__9,linha5_3__8,linha5_3__7,
              linha5_3__6,linha5_3__5,linha5_3__4,linha5_3__3,linha5_3__2,
              linha5_3__1,linha5_3__0}), .a1 ({linha6_2__63,linha6_2__62,
              linha6_2__61,linha6_2__60,linha6_2__59,linha6_2__58,linha6_2__57,
              linha6_2__56,linha6_2__55,linha6_2__54,linha6_2__53,linha6_2__52,
              linha6_2__51,linha6_2__50,linha6_2__49,linha6_2__48,linha6_2__47,
              linha6_2__46,linha6_2__45,linha6_2__44,linha6_2__43,linha6_2__42,
              linha6_2__41,linha6_2__40,linha6_2__39,linha6_2__38,linha6_2__37,
              linha6_2__36,linha6_2__35,linha6_2__34,linha6_2__33,linha6_2__32,
              linha6_2__31,linha6_2__30,linha6_2__29,linha6_2__28,linha6_2__27,
              linha6_2__26,linha6_2__25,linha6_2__24,linha6_2__23,linha6_2__22,
              linha6_2__21,linha6_2__20,linha6_2__19,linha6_2__18,linha6_2__17,
              linha6_2__16,linha6_2__15,linha6_2__14,linha6_2__13,linha6_2__12,
              linha6_2__11,linha6_2__10,linha6_2__9,linha6_2__8,linha6_2__7,
              linha6_2__6,linha6_2__5,linha6_2__4,linha6_2__3,linha6_2__2,
              linha6_2__1,linha6_2__0}), .a0 ({linha5_2__63,linha5_2__62,
              linha5_2__61,linha5_2__60,linha5_2__59,linha5_2__58,linha5_2__57,
              linha5_2__56,linha5_2__55,linha5_2__54,linha5_2__53,linha5_2__52,
              linha5_2__51,linha5_2__50,linha5_2__49,linha5_2__48,linha5_2__47,
              linha5_2__46,linha5_2__45,linha5_2__44,linha5_2__43,linha5_2__42,
              linha5_2__41,linha5_2__40,linha5_2__39,linha5_2__38,linha5_2__37,
              linha5_2__36,linha5_2__35,linha5_2__34,linha5_2__33,linha5_2__32,
              linha5_2__31,linha5_2__30,linha5_2__29,linha5_2__28,linha5_2__27,
              linha5_2__26,linha5_2__25,linha5_2__24,linha5_2__23,linha5_2__22,
              linha5_2__21,linha5_2__20,linha5_2__19,linha5_2__18,linha5_2__17,
              linha5_2__16,linha5_2__15,linha5_2__14,linha5_2__13,linha5_2__12,
              linha5_2__11,linha5_2__10,linha5_2__9,linha5_2__8,linha5_2__7,
              linha5_2__6,linha5_2__5,linha5_2__4,linha5_2__3,linha5_2__2,
              linha5_2__1,linha5_2__0}), .s (row_2_rowp_bni3_l)) ;
    Mux2x1_64 row_2_rowp_bni3_muxMin (.r ({linha6_3__63,linha6_3__62,
              linha6_3__61,linha6_3__60,linha6_3__59,linha6_3__58,linha6_3__57,
              linha6_3__56,linha6_3__55,linha6_3__54,linha6_3__53,linha6_3__52,
              linha6_3__51,linha6_3__50,linha6_3__49,linha6_3__48,linha6_3__47,
              linha6_3__46,linha6_3__45,linha6_3__44,linha6_3__43,linha6_3__42,
              linha6_3__41,linha6_3__40,linha6_3__39,linha6_3__38,linha6_3__37,
              linha6_3__36,linha6_3__35,linha6_3__34,linha6_3__33,linha6_3__32,
              linha6_3__31,linha6_3__30,linha6_3__29,linha6_3__28,linha6_3__27,
              linha6_3__26,linha6_3__25,linha6_3__24,linha6_3__23,linha6_3__22,
              linha6_3__21,linha6_3__20,linha6_3__19,linha6_3__18,linha6_3__17,
              linha6_3__16,linha6_3__15,linha6_3__14,linha6_3__13,linha6_3__12,
              linha6_3__11,linha6_3__10,linha6_3__9,linha6_3__8,linha6_3__7,
              linha6_3__6,linha6_3__5,linha6_3__4,linha6_3__3,linha6_3__2,
              linha6_3__1,linha6_3__0}), .a1 ({linha5_2__63,linha5_2__62,
              linha5_2__61,linha5_2__60,linha5_2__59,linha5_2__58,linha5_2__57,
              linha5_2__56,linha5_2__55,linha5_2__54,linha5_2__53,linha5_2__52,
              linha5_2__51,linha5_2__50,linha5_2__49,linha5_2__48,linha5_2__47,
              linha5_2__46,linha5_2__45,linha5_2__44,linha5_2__43,linha5_2__42,
              linha5_2__41,linha5_2__40,linha5_2__39,linha5_2__38,linha5_2__37,
              linha5_2__36,linha5_2__35,linha5_2__34,linha5_2__33,linha5_2__32,
              linha5_2__31,linha5_2__30,linha5_2__29,linha5_2__28,linha5_2__27,
              linha5_2__26,linha5_2__25,linha5_2__24,linha5_2__23,linha5_2__22,
              linha5_2__21,linha5_2__20,linha5_2__19,linha5_2__18,linha5_2__17,
              linha5_2__16,linha5_2__15,linha5_2__14,linha5_2__13,linha5_2__12,
              linha5_2__11,linha5_2__10,linha5_2__9,linha5_2__8,linha5_2__7,
              linha5_2__6,linha5_2__5,linha5_2__4,linha5_2__3,linha5_2__2,
              linha5_2__1,linha5_2__0}), .a0 ({linha6_2__63,linha6_2__62,
              linha6_2__61,linha6_2__60,linha6_2__59,linha6_2__58,linha6_2__57,
              linha6_2__56,linha6_2__55,linha6_2__54,linha6_2__53,linha6_2__52,
              linha6_2__51,linha6_2__50,linha6_2__49,linha6_2__48,linha6_2__47,
              linha6_2__46,linha6_2__45,linha6_2__44,linha6_2__43,linha6_2__42,
              linha6_2__41,linha6_2__40,linha6_2__39,linha6_2__38,linha6_2__37,
              linha6_2__36,linha6_2__35,linha6_2__34,linha6_2__33,linha6_2__32,
              linha6_2__31,linha6_2__30,linha6_2__29,linha6_2__28,linha6_2__27,
              linha6_2__26,linha6_2__25,linha6_2__24,linha6_2__23,linha6_2__22,
              linha6_2__21,linha6_2__20,linha6_2__19,linha6_2__18,linha6_2__17,
              linha6_2__16,linha6_2__15,linha6_2__14,linha6_2__13,linha6_2__12,
              linha6_2__11,linha6_2__10,linha6_2__9,linha6_2__8,linha6_2__7,
              linha6_2__6,linha6_2__5,linha6_2__4,linha6_2__3,linha6_2__2,
              linha6_2__1,linha6_2__0}), .s (row_2_rowp_bni3_l)) ;
    juntarComparadores_64 row_2_rowp_bni4_Comp (.g (\$dummy [10]), .l (
                          row_2_rowp_bni4_l), .a ({linha7_2__63,linha7_2__62,
                          linha7_2__61,linha7_2__60,linha7_2__59,linha7_2__58,
                          linha7_2__57,linha7_2__56,linha7_2__55,linha7_2__54,
                          linha7_2__53,linha7_2__52,linha7_2__51,linha7_2__50,
                          linha7_2__49,linha7_2__48,linha7_2__47,linha7_2__46,
                          linha7_2__45,linha7_2__44,linha7_2__43,linha7_2__42,
                          linha7_2__41,linha7_2__40,linha7_2__39,linha7_2__38,
                          linha7_2__37,linha7_2__36,linha7_2__35,linha7_2__34,
                          linha7_2__33,linha7_2__32,linha7_2__31,linha7_2__30,
                          linha7_2__29,linha7_2__28,linha7_2__27,linha7_2__26,
                          linha7_2__25,linha7_2__24,linha7_2__23,linha7_2__22,
                          linha7_2__21,linha7_2__20,linha7_2__19,linha7_2__18,
                          linha7_2__17,linha7_2__16,linha7_2__15,linha7_2__14,
                          linha7_2__13,linha7_2__12,linha7_2__11,linha7_2__10,
                          linha7_2__9,linha7_2__8,linha7_2__7,linha7_2__6,
                          linha7_2__5,linha7_2__4,linha7_2__3,linha7_2__2,
                          linha7_2__1,linha7_2__0}), .b ({linha8_1__63,
                          linha8_1__62,linha8_1__61,linha8_1__60,linha8_1__59,
                          linha8_1__58,linha8_1__57,linha8_1__56,linha8_1__55,
                          linha8_1__54,linha8_1__53,linha8_1__52,linha8_1__51,
                          linha8_1__50,linha8_1__49,linha8_1__48,linha8_1__47,
                          linha8_1__46,linha8_1__45,linha8_1__44,linha8_1__43,
                          linha8_1__42,linha8_1__41,linha8_1__40,linha8_1__39,
                          linha8_1__38,linha8_1__37,linha8_1__36,linha8_1__35,
                          linha8_1__34,linha8_1__33,linha8_1__32,linha8_1__31,
                          linha8_1__30,linha8_1__29,linha8_1__28,linha8_1__27,
                          linha8_1__26,linha8_1__25,linha8_1__24,linha8_1__23,
                          linha8_1__22,linha8_1__21,linha8_1__20,linha8_1__19,
                          linha8_1__18,linha8_1__17,linha8_1__16,linha8_1__15,
                          linha8_1__14,linha8_1__13,linha8_1__12,linha8_1__11,
                          linha8_1__10,linha8_1__9,linha8_1__8,linha8_1__7,
                          linha8_1__6,linha8_1__5,linha8_1__4,linha8_1__3,
                          linha8_1__2,linha8_1__1,linha8_1__0})) ;
    Mux2x1_64 row_2_rowp_bni4_muxMax (.r ({linha7_3__63,linha7_3__62,
              linha7_3__61,linha7_3__60,linha7_3__59,linha7_3__58,linha7_3__57,
              linha7_3__56,linha7_3__55,linha7_3__54,linha7_3__53,linha7_3__52,
              linha7_3__51,linha7_3__50,linha7_3__49,linha7_3__48,linha7_3__47,
              linha7_3__46,linha7_3__45,linha7_3__44,linha7_3__43,linha7_3__42,
              linha7_3__41,linha7_3__40,linha7_3__39,linha7_3__38,linha7_3__37,
              linha7_3__36,linha7_3__35,linha7_3__34,linha7_3__33,linha7_3__32,
              linha7_3__31,linha7_3__30,linha7_3__29,linha7_3__28,linha7_3__27,
              linha7_3__26,linha7_3__25,linha7_3__24,linha7_3__23,linha7_3__22,
              linha7_3__21,linha7_3__20,linha7_3__19,linha7_3__18,linha7_3__17,
              linha7_3__16,linha7_3__15,linha7_3__14,linha7_3__13,linha7_3__12,
              linha7_3__11,linha7_3__10,linha7_3__9,linha7_3__8,linha7_3__7,
              linha7_3__6,linha7_3__5,linha7_3__4,linha7_3__3,linha7_3__2,
              linha7_3__1,linha7_3__0}), .a1 ({linha8_1__63,linha8_1__62,
              linha8_1__61,linha8_1__60,linha8_1__59,linha8_1__58,linha8_1__57,
              linha8_1__56,linha8_1__55,linha8_1__54,linha8_1__53,linha8_1__52,
              linha8_1__51,linha8_1__50,linha8_1__49,linha8_1__48,linha8_1__47,
              linha8_1__46,linha8_1__45,linha8_1__44,linha8_1__43,linha8_1__42,
              linha8_1__41,linha8_1__40,linha8_1__39,linha8_1__38,linha8_1__37,
              linha8_1__36,linha8_1__35,linha8_1__34,linha8_1__33,linha8_1__32,
              linha8_1__31,linha8_1__30,linha8_1__29,linha8_1__28,linha8_1__27,
              linha8_1__26,linha8_1__25,linha8_1__24,linha8_1__23,linha8_1__22,
              linha8_1__21,linha8_1__20,linha8_1__19,linha8_1__18,linha8_1__17,
              linha8_1__16,linha8_1__15,linha8_1__14,linha8_1__13,linha8_1__12,
              linha8_1__11,linha8_1__10,linha8_1__9,linha8_1__8,linha8_1__7,
              linha8_1__6,linha8_1__5,linha8_1__4,linha8_1__3,linha8_1__2,
              linha8_1__1,linha8_1__0}), .a0 ({linha7_2__63,linha7_2__62,
              linha7_2__61,linha7_2__60,linha7_2__59,linha7_2__58,linha7_2__57,
              linha7_2__56,linha7_2__55,linha7_2__54,linha7_2__53,linha7_2__52,
              linha7_2__51,linha7_2__50,linha7_2__49,linha7_2__48,linha7_2__47,
              linha7_2__46,linha7_2__45,linha7_2__44,linha7_2__43,linha7_2__42,
              linha7_2__41,linha7_2__40,linha7_2__39,linha7_2__38,linha7_2__37,
              linha7_2__36,linha7_2__35,linha7_2__34,linha7_2__33,linha7_2__32,
              linha7_2__31,linha7_2__30,linha7_2__29,linha7_2__28,linha7_2__27,
              linha7_2__26,linha7_2__25,linha7_2__24,linha7_2__23,linha7_2__22,
              linha7_2__21,linha7_2__20,linha7_2__19,linha7_2__18,linha7_2__17,
              linha7_2__16,linha7_2__15,linha7_2__14,linha7_2__13,linha7_2__12,
              linha7_2__11,linha7_2__10,linha7_2__9,linha7_2__8,linha7_2__7,
              linha7_2__6,linha7_2__5,linha7_2__4,linha7_2__3,linha7_2__2,
              linha7_2__1,linha7_2__0}), .s (row_2_rowp_bni4_l)) ;
    Mux2x1_64 row_2_rowp_bni4_muxMin (.r ({linha8_2__63,linha8_2__62,
              linha8_2__61,linha8_2__60,linha8_2__59,linha8_2__58,linha8_2__57,
              linha8_2__56,linha8_2__55,linha8_2__54,linha8_2__53,linha8_2__52,
              linha8_2__51,linha8_2__50,linha8_2__49,linha8_2__48,linha8_2__47,
              linha8_2__46,linha8_2__45,linha8_2__44,linha8_2__43,linha8_2__42,
              linha8_2__41,linha8_2__40,linha8_2__39,linha8_2__38,linha8_2__37,
              linha8_2__36,linha8_2__35,linha8_2__34,linha8_2__33,linha8_2__32,
              linha8_2__31,linha8_2__30,linha8_2__29,linha8_2__28,linha8_2__27,
              linha8_2__26,linha8_2__25,linha8_2__24,linha8_2__23,linha8_2__22,
              linha8_2__21,linha8_2__20,linha8_2__19,linha8_2__18,linha8_2__17,
              linha8_2__16,linha8_2__15,linha8_2__14,linha8_2__13,linha8_2__12,
              linha8_2__11,linha8_2__10,linha8_2__9,linha8_2__8,linha8_2__7,
              linha8_2__6,linha8_2__5,linha8_2__4,linha8_2__3,linha8_2__2,
              linha8_2__1,linha8_2__0}), .a1 ({linha7_2__63,linha7_2__62,
              linha7_2__61,linha7_2__60,linha7_2__59,linha7_2__58,linha7_2__57,
              linha7_2__56,linha7_2__55,linha7_2__54,linha7_2__53,linha7_2__52,
              linha7_2__51,linha7_2__50,linha7_2__49,linha7_2__48,linha7_2__47,
              linha7_2__46,linha7_2__45,linha7_2__44,linha7_2__43,linha7_2__42,
              linha7_2__41,linha7_2__40,linha7_2__39,linha7_2__38,linha7_2__37,
              linha7_2__36,linha7_2__35,linha7_2__34,linha7_2__33,linha7_2__32,
              linha7_2__31,linha7_2__30,linha7_2__29,linha7_2__28,linha7_2__27,
              linha7_2__26,linha7_2__25,linha7_2__24,linha7_2__23,linha7_2__22,
              linha7_2__21,linha7_2__20,linha7_2__19,linha7_2__18,linha7_2__17,
              linha7_2__16,linha7_2__15,linha7_2__14,linha7_2__13,linha7_2__12,
              linha7_2__11,linha7_2__10,linha7_2__9,linha7_2__8,linha7_2__7,
              linha7_2__6,linha7_2__5,linha7_2__4,linha7_2__3,linha7_2__2,
              linha7_2__1,linha7_2__0}), .a0 ({linha8_1__63,linha8_1__62,
              linha8_1__61,linha8_1__60,linha8_1__59,linha8_1__58,linha8_1__57,
              linha8_1__56,linha8_1__55,linha8_1__54,linha8_1__53,linha8_1__52,
              linha8_1__51,linha8_1__50,linha8_1__49,linha8_1__48,linha8_1__47,
              linha8_1__46,linha8_1__45,linha8_1__44,linha8_1__43,linha8_1__42,
              linha8_1__41,linha8_1__40,linha8_1__39,linha8_1__38,linha8_1__37,
              linha8_1__36,linha8_1__35,linha8_1__34,linha8_1__33,linha8_1__32,
              linha8_1__31,linha8_1__30,linha8_1__29,linha8_1__28,linha8_1__27,
              linha8_1__26,linha8_1__25,linha8_1__24,linha8_1__23,linha8_1__22,
              linha8_1__21,linha8_1__20,linha8_1__19,linha8_1__18,linha8_1__17,
              linha8_1__16,linha8_1__15,linha8_1__14,linha8_1__13,linha8_1__12,
              linha8_1__11,linha8_1__10,linha8_1__9,linha8_1__8,linha8_1__7,
              linha8_1__6,linha8_1__5,linha8_1__4,linha8_1__3,linha8_1__2,
              linha8_1__1,linha8_1__0}), .s (row_2_rowp_bni4_l)) ;
    juntarComparadores_64 row_3_rowi_bni1_Comp (.g (\$dummy [11]), .l (
                          row_3_rowi_bni1_l), .a ({linha2_3__63,linha2_3__62,
                          linha2_3__61,linha2_3__60,linha2_3__59,linha2_3__58,
                          linha2_3__57,linha2_3__56,linha2_3__55,linha2_3__54,
                          linha2_3__53,linha2_3__52,linha2_3__51,linha2_3__50,
                          linha2_3__49,linha2_3__48,linha2_3__47,linha2_3__46,
                          linha2_3__45,linha2_3__44,linha2_3__43,linha2_3__42,
                          linha2_3__41,linha2_3__40,linha2_3__39,linha2_3__38,
                          linha2_3__37,linha2_3__36,linha2_3__35,linha2_3__34,
                          linha2_3__33,linha2_3__32,linha2_3__31,linha2_3__30,
                          linha2_3__29,linha2_3__28,linha2_3__27,linha2_3__26,
                          linha2_3__25,linha2_3__24,linha2_3__23,linha2_3__22,
                          linha2_3__21,linha2_3__20,linha2_3__19,linha2_3__18,
                          linha2_3__17,linha2_3__16,linha2_3__15,linha2_3__14,
                          linha2_3__13,linha2_3__12,linha2_3__11,linha2_3__10,
                          linha2_3__9,linha2_3__8,linha2_3__7,linha2_3__6,
                          linha2_3__5,linha2_3__4,linha2_3__3,linha2_3__2,
                          linha2_3__1,linha2_3__0}), .b ({linha3_3__63,
                          linha3_3__62,linha3_3__61,linha3_3__60,linha3_3__59,
                          linha3_3__58,linha3_3__57,linha3_3__56,linha3_3__55,
                          linha3_3__54,linha3_3__53,linha3_3__52,linha3_3__51,
                          linha3_3__50,linha3_3__49,linha3_3__48,linha3_3__47,
                          linha3_3__46,linha3_3__45,linha3_3__44,linha3_3__43,
                          linha3_3__42,linha3_3__41,linha3_3__40,linha3_3__39,
                          linha3_3__38,linha3_3__37,linha3_3__36,linha3_3__35,
                          linha3_3__34,linha3_3__33,linha3_3__32,linha3_3__31,
                          linha3_3__30,linha3_3__29,linha3_3__28,linha3_3__27,
                          linha3_3__26,linha3_3__25,linha3_3__24,linha3_3__23,
                          linha3_3__22,linha3_3__21,linha3_3__20,linha3_3__19,
                          linha3_3__18,linha3_3__17,linha3_3__16,linha3_3__15,
                          linha3_3__14,linha3_3__13,linha3_3__12,linha3_3__11,
                          linha3_3__10,linha3_3__9,linha3_3__8,linha3_3__7,
                          linha3_3__6,linha3_3__5,linha3_3__4,linha3_3__3,
                          linha3_3__2,linha3_3__1,linha3_3__0})) ;
    Mux2x1_64 row_3_rowi_bni1_muxMax (.r ({linha2_4__63,linha2_4__62,
              linha2_4__61,linha2_4__60,linha2_4__59,linha2_4__58,linha2_4__57,
              linha2_4__56,linha2_4__55,linha2_4__54,linha2_4__53,linha2_4__52,
              linha2_4__51,linha2_4__50,linha2_4__49,linha2_4__48,linha2_4__47,
              linha2_4__46,linha2_4__45,linha2_4__44,linha2_4__43,linha2_4__42,
              linha2_4__41,linha2_4__40,linha2_4__39,linha2_4__38,linha2_4__37,
              linha2_4__36,linha2_4__35,linha2_4__34,linha2_4__33,linha2_4__32,
              linha2_4__31,linha2_4__30,linha2_4__29,linha2_4__28,linha2_4__27,
              linha2_4__26,linha2_4__25,linha2_4__24,linha2_4__23,linha2_4__22,
              linha2_4__21,linha2_4__20,linha2_4__19,linha2_4__18,linha2_4__17,
              linha2_4__16,linha2_4__15,linha2_4__14,linha2_4__13,linha2_4__12,
              linha2_4__11,linha2_4__10,linha2_4__9,linha2_4__8,linha2_4__7,
              linha2_4__6,linha2_4__5,linha2_4__4,linha2_4__3,linha2_4__2,
              linha2_4__1,linha2_4__0}), .a1 ({linha3_3__63,linha3_3__62,
              linha3_3__61,linha3_3__60,linha3_3__59,linha3_3__58,linha3_3__57,
              linha3_3__56,linha3_3__55,linha3_3__54,linha3_3__53,linha3_3__52,
              linha3_3__51,linha3_3__50,linha3_3__49,linha3_3__48,linha3_3__47,
              linha3_3__46,linha3_3__45,linha3_3__44,linha3_3__43,linha3_3__42,
              linha3_3__41,linha3_3__40,linha3_3__39,linha3_3__38,linha3_3__37,
              linha3_3__36,linha3_3__35,linha3_3__34,linha3_3__33,linha3_3__32,
              linha3_3__31,linha3_3__30,linha3_3__29,linha3_3__28,linha3_3__27,
              linha3_3__26,linha3_3__25,linha3_3__24,linha3_3__23,linha3_3__22,
              linha3_3__21,linha3_3__20,linha3_3__19,linha3_3__18,linha3_3__17,
              linha3_3__16,linha3_3__15,linha3_3__14,linha3_3__13,linha3_3__12,
              linha3_3__11,linha3_3__10,linha3_3__9,linha3_3__8,linha3_3__7,
              linha3_3__6,linha3_3__5,linha3_3__4,linha3_3__3,linha3_3__2,
              linha3_3__1,linha3_3__0}), .a0 ({linha2_3__63,linha2_3__62,
              linha2_3__61,linha2_3__60,linha2_3__59,linha2_3__58,linha2_3__57,
              linha2_3__56,linha2_3__55,linha2_3__54,linha2_3__53,linha2_3__52,
              linha2_3__51,linha2_3__50,linha2_3__49,linha2_3__48,linha2_3__47,
              linha2_3__46,linha2_3__45,linha2_3__44,linha2_3__43,linha2_3__42,
              linha2_3__41,linha2_3__40,linha2_3__39,linha2_3__38,linha2_3__37,
              linha2_3__36,linha2_3__35,linha2_3__34,linha2_3__33,linha2_3__32,
              linha2_3__31,linha2_3__30,linha2_3__29,linha2_3__28,linha2_3__27,
              linha2_3__26,linha2_3__25,linha2_3__24,linha2_3__23,linha2_3__22,
              linha2_3__21,linha2_3__20,linha2_3__19,linha2_3__18,linha2_3__17,
              linha2_3__16,linha2_3__15,linha2_3__14,linha2_3__13,linha2_3__12,
              linha2_3__11,linha2_3__10,linha2_3__9,linha2_3__8,linha2_3__7,
              linha2_3__6,linha2_3__5,linha2_3__4,linha2_3__3,linha2_3__2,
              linha2_3__1,linha2_3__0}), .s (row_3_rowi_bni1_l)) ;
    Mux2x1_64 row_3_rowi_bni1_muxMin (.r ({linha3_4__63,linha3_4__62,
              linha3_4__61,linha3_4__60,linha3_4__59,linha3_4__58,linha3_4__57,
              linha3_4__56,linha3_4__55,linha3_4__54,linha3_4__53,linha3_4__52,
              linha3_4__51,linha3_4__50,linha3_4__49,linha3_4__48,linha3_4__47,
              linha3_4__46,linha3_4__45,linha3_4__44,linha3_4__43,linha3_4__42,
              linha3_4__41,linha3_4__40,linha3_4__39,linha3_4__38,linha3_4__37,
              linha3_4__36,linha3_4__35,linha3_4__34,linha3_4__33,linha3_4__32,
              linha3_4__31,linha3_4__30,linha3_4__29,linha3_4__28,linha3_4__27,
              linha3_4__26,linha3_4__25,linha3_4__24,linha3_4__23,linha3_4__22,
              linha3_4__21,linha3_4__20,linha3_4__19,linha3_4__18,linha3_4__17,
              linha3_4__16,linha3_4__15,linha3_4__14,linha3_4__13,linha3_4__12,
              linha3_4__11,linha3_4__10,linha3_4__9,linha3_4__8,linha3_4__7,
              linha3_4__6,linha3_4__5,linha3_4__4,linha3_4__3,linha3_4__2,
              linha3_4__1,linha3_4__0}), .a1 ({linha2_3__63,linha2_3__62,
              linha2_3__61,linha2_3__60,linha2_3__59,linha2_3__58,linha2_3__57,
              linha2_3__56,linha2_3__55,linha2_3__54,linha2_3__53,linha2_3__52,
              linha2_3__51,linha2_3__50,linha2_3__49,linha2_3__48,linha2_3__47,
              linha2_3__46,linha2_3__45,linha2_3__44,linha2_3__43,linha2_3__42,
              linha2_3__41,linha2_3__40,linha2_3__39,linha2_3__38,linha2_3__37,
              linha2_3__36,linha2_3__35,linha2_3__34,linha2_3__33,linha2_3__32,
              linha2_3__31,linha2_3__30,linha2_3__29,linha2_3__28,linha2_3__27,
              linha2_3__26,linha2_3__25,linha2_3__24,linha2_3__23,linha2_3__22,
              linha2_3__21,linha2_3__20,linha2_3__19,linha2_3__18,linha2_3__17,
              linha2_3__16,linha2_3__15,linha2_3__14,linha2_3__13,linha2_3__12,
              linha2_3__11,linha2_3__10,linha2_3__9,linha2_3__8,linha2_3__7,
              linha2_3__6,linha2_3__5,linha2_3__4,linha2_3__3,linha2_3__2,
              linha2_3__1,linha2_3__0}), .a0 ({linha3_3__63,linha3_3__62,
              linha3_3__61,linha3_3__60,linha3_3__59,linha3_3__58,linha3_3__57,
              linha3_3__56,linha3_3__55,linha3_3__54,linha3_3__53,linha3_3__52,
              linha3_3__51,linha3_3__50,linha3_3__49,linha3_3__48,linha3_3__47,
              linha3_3__46,linha3_3__45,linha3_3__44,linha3_3__43,linha3_3__42,
              linha3_3__41,linha3_3__40,linha3_3__39,linha3_3__38,linha3_3__37,
              linha3_3__36,linha3_3__35,linha3_3__34,linha3_3__33,linha3_3__32,
              linha3_3__31,linha3_3__30,linha3_3__29,linha3_3__28,linha3_3__27,
              linha3_3__26,linha3_3__25,linha3_3__24,linha3_3__23,linha3_3__22,
              linha3_3__21,linha3_3__20,linha3_3__19,linha3_3__18,linha3_3__17,
              linha3_3__16,linha3_3__15,linha3_3__14,linha3_3__13,linha3_3__12,
              linha3_3__11,linha3_3__10,linha3_3__9,linha3_3__8,linha3_3__7,
              linha3_3__6,linha3_3__5,linha3_3__4,linha3_3__3,linha3_3__2,
              linha3_3__1,linha3_3__0}), .s (row_3_rowi_bni1_l)) ;
    juntarComparadores_64 row_3_rowi_bni2_Comp (.g (\$dummy [12]), .l (
                          row_3_rowi_bni2_l), .a ({linha4_3__63,linha4_3__62,
                          linha4_3__61,linha4_3__60,linha4_3__59,linha4_3__58,
                          linha4_3__57,linha4_3__56,linha4_3__55,linha4_3__54,
                          linha4_3__53,linha4_3__52,linha4_3__51,linha4_3__50,
                          linha4_3__49,linha4_3__48,linha4_3__47,linha4_3__46,
                          linha4_3__45,linha4_3__44,linha4_3__43,linha4_3__42,
                          linha4_3__41,linha4_3__40,linha4_3__39,linha4_3__38,
                          linha4_3__37,linha4_3__36,linha4_3__35,linha4_3__34,
                          linha4_3__33,linha4_3__32,linha4_3__31,linha4_3__30,
                          linha4_3__29,linha4_3__28,linha4_3__27,linha4_3__26,
                          linha4_3__25,linha4_3__24,linha4_3__23,linha4_3__22,
                          linha4_3__21,linha4_3__20,linha4_3__19,linha4_3__18,
                          linha4_3__17,linha4_3__16,linha4_3__15,linha4_3__14,
                          linha4_3__13,linha4_3__12,linha4_3__11,linha4_3__10,
                          linha4_3__9,linha4_3__8,linha4_3__7,linha4_3__6,
                          linha4_3__5,linha4_3__4,linha4_3__3,linha4_3__2,
                          linha4_3__1,linha4_3__0}), .b ({linha5_3__63,
                          linha5_3__62,linha5_3__61,linha5_3__60,linha5_3__59,
                          linha5_3__58,linha5_3__57,linha5_3__56,linha5_3__55,
                          linha5_3__54,linha5_3__53,linha5_3__52,linha5_3__51,
                          linha5_3__50,linha5_3__49,linha5_3__48,linha5_3__47,
                          linha5_3__46,linha5_3__45,linha5_3__44,linha5_3__43,
                          linha5_3__42,linha5_3__41,linha5_3__40,linha5_3__39,
                          linha5_3__38,linha5_3__37,linha5_3__36,linha5_3__35,
                          linha5_3__34,linha5_3__33,linha5_3__32,linha5_3__31,
                          linha5_3__30,linha5_3__29,linha5_3__28,linha5_3__27,
                          linha5_3__26,linha5_3__25,linha5_3__24,linha5_3__23,
                          linha5_3__22,linha5_3__21,linha5_3__20,linha5_3__19,
                          linha5_3__18,linha5_3__17,linha5_3__16,linha5_3__15,
                          linha5_3__14,linha5_3__13,linha5_3__12,linha5_3__11,
                          linha5_3__10,linha5_3__9,linha5_3__8,linha5_3__7,
                          linha5_3__6,linha5_3__5,linha5_3__4,linha5_3__3,
                          linha5_3__2,linha5_3__1,linha5_3__0})) ;
    Mux2x1_64 row_3_rowi_bni2_muxMax (.r ({linha4_4__63,linha4_4__62,
              linha4_4__61,linha4_4__60,linha4_4__59,linha4_4__58,linha4_4__57,
              linha4_4__56,linha4_4__55,linha4_4__54,linha4_4__53,linha4_4__52,
              linha4_4__51,linha4_4__50,linha4_4__49,linha4_4__48,linha4_4__47,
              linha4_4__46,linha4_4__45,linha4_4__44,linha4_4__43,linha4_4__42,
              linha4_4__41,linha4_4__40,linha4_4__39,linha4_4__38,linha4_4__37,
              linha4_4__36,linha4_4__35,linha4_4__34,linha4_4__33,linha4_4__32,
              linha4_4__31,linha4_4__30,linha4_4__29,linha4_4__28,linha4_4__27,
              linha4_4__26,linha4_4__25,linha4_4__24,linha4_4__23,linha4_4__22,
              linha4_4__21,linha4_4__20,linha4_4__19,linha4_4__18,linha4_4__17,
              linha4_4__16,linha4_4__15,linha4_4__14,linha4_4__13,linha4_4__12,
              linha4_4__11,linha4_4__10,linha4_4__9,linha4_4__8,linha4_4__7,
              linha4_4__6,linha4_4__5,linha4_4__4,linha4_4__3,linha4_4__2,
              linha4_4__1,linha4_4__0}), .a1 ({linha5_3__63,linha5_3__62,
              linha5_3__61,linha5_3__60,linha5_3__59,linha5_3__58,linha5_3__57,
              linha5_3__56,linha5_3__55,linha5_3__54,linha5_3__53,linha5_3__52,
              linha5_3__51,linha5_3__50,linha5_3__49,linha5_3__48,linha5_3__47,
              linha5_3__46,linha5_3__45,linha5_3__44,linha5_3__43,linha5_3__42,
              linha5_3__41,linha5_3__40,linha5_3__39,linha5_3__38,linha5_3__37,
              linha5_3__36,linha5_3__35,linha5_3__34,linha5_3__33,linha5_3__32,
              linha5_3__31,linha5_3__30,linha5_3__29,linha5_3__28,linha5_3__27,
              linha5_3__26,linha5_3__25,linha5_3__24,linha5_3__23,linha5_3__22,
              linha5_3__21,linha5_3__20,linha5_3__19,linha5_3__18,linha5_3__17,
              linha5_3__16,linha5_3__15,linha5_3__14,linha5_3__13,linha5_3__12,
              linha5_3__11,linha5_3__10,linha5_3__9,linha5_3__8,linha5_3__7,
              linha5_3__6,linha5_3__5,linha5_3__4,linha5_3__3,linha5_3__2,
              linha5_3__1,linha5_3__0}), .a0 ({linha4_3__63,linha4_3__62,
              linha4_3__61,linha4_3__60,linha4_3__59,linha4_3__58,linha4_3__57,
              linha4_3__56,linha4_3__55,linha4_3__54,linha4_3__53,linha4_3__52,
              linha4_3__51,linha4_3__50,linha4_3__49,linha4_3__48,linha4_3__47,
              linha4_3__46,linha4_3__45,linha4_3__44,linha4_3__43,linha4_3__42,
              linha4_3__41,linha4_3__40,linha4_3__39,linha4_3__38,linha4_3__37,
              linha4_3__36,linha4_3__35,linha4_3__34,linha4_3__33,linha4_3__32,
              linha4_3__31,linha4_3__30,linha4_3__29,linha4_3__28,linha4_3__27,
              linha4_3__26,linha4_3__25,linha4_3__24,linha4_3__23,linha4_3__22,
              linha4_3__21,linha4_3__20,linha4_3__19,linha4_3__18,linha4_3__17,
              linha4_3__16,linha4_3__15,linha4_3__14,linha4_3__13,linha4_3__12,
              linha4_3__11,linha4_3__10,linha4_3__9,linha4_3__8,linha4_3__7,
              linha4_3__6,linha4_3__5,linha4_3__4,linha4_3__3,linha4_3__2,
              linha4_3__1,linha4_3__0}), .s (row_3_rowi_bni2_l)) ;
    Mux2x1_64 row_3_rowi_bni2_muxMin (.r ({linha5_4__63,linha5_4__62,
              linha5_4__61,linha5_4__60,linha5_4__59,linha5_4__58,linha5_4__57,
              linha5_4__56,linha5_4__55,linha5_4__54,linha5_4__53,linha5_4__52,
              linha5_4__51,linha5_4__50,linha5_4__49,linha5_4__48,linha5_4__47,
              linha5_4__46,linha5_4__45,linha5_4__44,linha5_4__43,linha5_4__42,
              linha5_4__41,linha5_4__40,linha5_4__39,linha5_4__38,linha5_4__37,
              linha5_4__36,linha5_4__35,linha5_4__34,linha5_4__33,linha5_4__32,
              linha5_4__31,linha5_4__30,linha5_4__29,linha5_4__28,linha5_4__27,
              linha5_4__26,linha5_4__25,linha5_4__24,linha5_4__23,linha5_4__22,
              linha5_4__21,linha5_4__20,linha5_4__19,linha5_4__18,linha5_4__17,
              linha5_4__16,linha5_4__15,linha5_4__14,linha5_4__13,linha5_4__12,
              linha5_4__11,linha5_4__10,linha5_4__9,linha5_4__8,linha5_4__7,
              linha5_4__6,linha5_4__5,linha5_4__4,linha5_4__3,linha5_4__2,
              linha5_4__1,linha5_4__0}), .a1 ({linha4_3__63,linha4_3__62,
              linha4_3__61,linha4_3__60,linha4_3__59,linha4_3__58,linha4_3__57,
              linha4_3__56,linha4_3__55,linha4_3__54,linha4_3__53,linha4_3__52,
              linha4_3__51,linha4_3__50,linha4_3__49,linha4_3__48,linha4_3__47,
              linha4_3__46,linha4_3__45,linha4_3__44,linha4_3__43,linha4_3__42,
              linha4_3__41,linha4_3__40,linha4_3__39,linha4_3__38,linha4_3__37,
              linha4_3__36,linha4_3__35,linha4_3__34,linha4_3__33,linha4_3__32,
              linha4_3__31,linha4_3__30,linha4_3__29,linha4_3__28,linha4_3__27,
              linha4_3__26,linha4_3__25,linha4_3__24,linha4_3__23,linha4_3__22,
              linha4_3__21,linha4_3__20,linha4_3__19,linha4_3__18,linha4_3__17,
              linha4_3__16,linha4_3__15,linha4_3__14,linha4_3__13,linha4_3__12,
              linha4_3__11,linha4_3__10,linha4_3__9,linha4_3__8,linha4_3__7,
              linha4_3__6,linha4_3__5,linha4_3__4,linha4_3__3,linha4_3__2,
              linha4_3__1,linha4_3__0}), .a0 ({linha5_3__63,linha5_3__62,
              linha5_3__61,linha5_3__60,linha5_3__59,linha5_3__58,linha5_3__57,
              linha5_3__56,linha5_3__55,linha5_3__54,linha5_3__53,linha5_3__52,
              linha5_3__51,linha5_3__50,linha5_3__49,linha5_3__48,linha5_3__47,
              linha5_3__46,linha5_3__45,linha5_3__44,linha5_3__43,linha5_3__42,
              linha5_3__41,linha5_3__40,linha5_3__39,linha5_3__38,linha5_3__37,
              linha5_3__36,linha5_3__35,linha5_3__34,linha5_3__33,linha5_3__32,
              linha5_3__31,linha5_3__30,linha5_3__29,linha5_3__28,linha5_3__27,
              linha5_3__26,linha5_3__25,linha5_3__24,linha5_3__23,linha5_3__22,
              linha5_3__21,linha5_3__20,linha5_3__19,linha5_3__18,linha5_3__17,
              linha5_3__16,linha5_3__15,linha5_3__14,linha5_3__13,linha5_3__12,
              linha5_3__11,linha5_3__10,linha5_3__9,linha5_3__8,linha5_3__7,
              linha5_3__6,linha5_3__5,linha5_3__4,linha5_3__3,linha5_3__2,
              linha5_3__1,linha5_3__0}), .s (row_3_rowi_bni2_l)) ;
    juntarComparadores_64 row_3_rowi_bni3_Comp (.g (\$dummy [13]), .l (
                          row_3_rowi_bni3_l), .a ({linha6_3__63,linha6_3__62,
                          linha6_3__61,linha6_3__60,linha6_3__59,linha6_3__58,
                          linha6_3__57,linha6_3__56,linha6_3__55,linha6_3__54,
                          linha6_3__53,linha6_3__52,linha6_3__51,linha6_3__50,
                          linha6_3__49,linha6_3__48,linha6_3__47,linha6_3__46,
                          linha6_3__45,linha6_3__44,linha6_3__43,linha6_3__42,
                          linha6_3__41,linha6_3__40,linha6_3__39,linha6_3__38,
                          linha6_3__37,linha6_3__36,linha6_3__35,linha6_3__34,
                          linha6_3__33,linha6_3__32,linha6_3__31,linha6_3__30,
                          linha6_3__29,linha6_3__28,linha6_3__27,linha6_3__26,
                          linha6_3__25,linha6_3__24,linha6_3__23,linha6_3__22,
                          linha6_3__21,linha6_3__20,linha6_3__19,linha6_3__18,
                          linha6_3__17,linha6_3__16,linha6_3__15,linha6_3__14,
                          linha6_3__13,linha6_3__12,linha6_3__11,linha6_3__10,
                          linha6_3__9,linha6_3__8,linha6_3__7,linha6_3__6,
                          linha6_3__5,linha6_3__4,linha6_3__3,linha6_3__2,
                          linha6_3__1,linha6_3__0}), .b ({linha7_3__63,
                          linha7_3__62,linha7_3__61,linha7_3__60,linha7_3__59,
                          linha7_3__58,linha7_3__57,linha7_3__56,linha7_3__55,
                          linha7_3__54,linha7_3__53,linha7_3__52,linha7_3__51,
                          linha7_3__50,linha7_3__49,linha7_3__48,linha7_3__47,
                          linha7_3__46,linha7_3__45,linha7_3__44,linha7_3__43,
                          linha7_3__42,linha7_3__41,linha7_3__40,linha7_3__39,
                          linha7_3__38,linha7_3__37,linha7_3__36,linha7_3__35,
                          linha7_3__34,linha7_3__33,linha7_3__32,linha7_3__31,
                          linha7_3__30,linha7_3__29,linha7_3__28,linha7_3__27,
                          linha7_3__26,linha7_3__25,linha7_3__24,linha7_3__23,
                          linha7_3__22,linha7_3__21,linha7_3__20,linha7_3__19,
                          linha7_3__18,linha7_3__17,linha7_3__16,linha7_3__15,
                          linha7_3__14,linha7_3__13,linha7_3__12,linha7_3__11,
                          linha7_3__10,linha7_3__9,linha7_3__8,linha7_3__7,
                          linha7_3__6,linha7_3__5,linha7_3__4,linha7_3__3,
                          linha7_3__2,linha7_3__1,linha7_3__0})) ;
    Mux2x1_64 row_3_rowi_bni3_muxMax (.r ({linha6_4__63,linha6_4__62,
              linha6_4__61,linha6_4__60,linha6_4__59,linha6_4__58,linha6_4__57,
              linha6_4__56,linha6_4__55,linha6_4__54,linha6_4__53,linha6_4__52,
              linha6_4__51,linha6_4__50,linha6_4__49,linha6_4__48,linha6_4__47,
              linha6_4__46,linha6_4__45,linha6_4__44,linha6_4__43,linha6_4__42,
              linha6_4__41,linha6_4__40,linha6_4__39,linha6_4__38,linha6_4__37,
              linha6_4__36,linha6_4__35,linha6_4__34,linha6_4__33,linha6_4__32,
              linha6_4__31,linha6_4__30,linha6_4__29,linha6_4__28,linha6_4__27,
              linha6_4__26,linha6_4__25,linha6_4__24,linha6_4__23,linha6_4__22,
              linha6_4__21,linha6_4__20,linha6_4__19,linha6_4__18,linha6_4__17,
              linha6_4__16,linha6_4__15,linha6_4__14,linha6_4__13,linha6_4__12,
              linha6_4__11,linha6_4__10,linha6_4__9,linha6_4__8,linha6_4__7,
              linha6_4__6,linha6_4__5,linha6_4__4,linha6_4__3,linha6_4__2,
              linha6_4__1,linha6_4__0}), .a1 ({linha7_3__63,linha7_3__62,
              linha7_3__61,linha7_3__60,linha7_3__59,linha7_3__58,linha7_3__57,
              linha7_3__56,linha7_3__55,linha7_3__54,linha7_3__53,linha7_3__52,
              linha7_3__51,linha7_3__50,linha7_3__49,linha7_3__48,linha7_3__47,
              linha7_3__46,linha7_3__45,linha7_3__44,linha7_3__43,linha7_3__42,
              linha7_3__41,linha7_3__40,linha7_3__39,linha7_3__38,linha7_3__37,
              linha7_3__36,linha7_3__35,linha7_3__34,linha7_3__33,linha7_3__32,
              linha7_3__31,linha7_3__30,linha7_3__29,linha7_3__28,linha7_3__27,
              linha7_3__26,linha7_3__25,linha7_3__24,linha7_3__23,linha7_3__22,
              linha7_3__21,linha7_3__20,linha7_3__19,linha7_3__18,linha7_3__17,
              linha7_3__16,linha7_3__15,linha7_3__14,linha7_3__13,linha7_3__12,
              linha7_3__11,linha7_3__10,linha7_3__9,linha7_3__8,linha7_3__7,
              linha7_3__6,linha7_3__5,linha7_3__4,linha7_3__3,linha7_3__2,
              linha7_3__1,linha7_3__0}), .a0 ({linha6_3__63,linha6_3__62,
              linha6_3__61,linha6_3__60,linha6_3__59,linha6_3__58,linha6_3__57,
              linha6_3__56,linha6_3__55,linha6_3__54,linha6_3__53,linha6_3__52,
              linha6_3__51,linha6_3__50,linha6_3__49,linha6_3__48,linha6_3__47,
              linha6_3__46,linha6_3__45,linha6_3__44,linha6_3__43,linha6_3__42,
              linha6_3__41,linha6_3__40,linha6_3__39,linha6_3__38,linha6_3__37,
              linha6_3__36,linha6_3__35,linha6_3__34,linha6_3__33,linha6_3__32,
              linha6_3__31,linha6_3__30,linha6_3__29,linha6_3__28,linha6_3__27,
              linha6_3__26,linha6_3__25,linha6_3__24,linha6_3__23,linha6_3__22,
              linha6_3__21,linha6_3__20,linha6_3__19,linha6_3__18,linha6_3__17,
              linha6_3__16,linha6_3__15,linha6_3__14,linha6_3__13,linha6_3__12,
              linha6_3__11,linha6_3__10,linha6_3__9,linha6_3__8,linha6_3__7,
              linha6_3__6,linha6_3__5,linha6_3__4,linha6_3__3,linha6_3__2,
              linha6_3__1,linha6_3__0}), .s (row_3_rowi_bni3_l)) ;
    Mux2x1_64 row_3_rowi_bni3_muxMin (.r ({linha7_4__63,linha7_4__62,
              linha7_4__61,linha7_4__60,linha7_4__59,linha7_4__58,linha7_4__57,
              linha7_4__56,linha7_4__55,linha7_4__54,linha7_4__53,linha7_4__52,
              linha7_4__51,linha7_4__50,linha7_4__49,linha7_4__48,linha7_4__47,
              linha7_4__46,linha7_4__45,linha7_4__44,linha7_4__43,linha7_4__42,
              linha7_4__41,linha7_4__40,linha7_4__39,linha7_4__38,linha7_4__37,
              linha7_4__36,linha7_4__35,linha7_4__34,linha7_4__33,linha7_4__32,
              linha7_4__31,linha7_4__30,linha7_4__29,linha7_4__28,linha7_4__27,
              linha7_4__26,linha7_4__25,linha7_4__24,linha7_4__23,linha7_4__22,
              linha7_4__21,linha7_4__20,linha7_4__19,linha7_4__18,linha7_4__17,
              linha7_4__16,linha7_4__15,linha7_4__14,linha7_4__13,linha7_4__12,
              linha7_4__11,linha7_4__10,linha7_4__9,linha7_4__8,linha7_4__7,
              linha7_4__6,linha7_4__5,linha7_4__4,linha7_4__3,linha7_4__2,
              linha7_4__1,linha7_4__0}), .a1 ({linha6_3__63,linha6_3__62,
              linha6_3__61,linha6_3__60,linha6_3__59,linha6_3__58,linha6_3__57,
              linha6_3__56,linha6_3__55,linha6_3__54,linha6_3__53,linha6_3__52,
              linha6_3__51,linha6_3__50,linha6_3__49,linha6_3__48,linha6_3__47,
              linha6_3__46,linha6_3__45,linha6_3__44,linha6_3__43,linha6_3__42,
              linha6_3__41,linha6_3__40,linha6_3__39,linha6_3__38,linha6_3__37,
              linha6_3__36,linha6_3__35,linha6_3__34,linha6_3__33,linha6_3__32,
              linha6_3__31,linha6_3__30,linha6_3__29,linha6_3__28,linha6_3__27,
              linha6_3__26,linha6_3__25,linha6_3__24,linha6_3__23,linha6_3__22,
              linha6_3__21,linha6_3__20,linha6_3__19,linha6_3__18,linha6_3__17,
              linha6_3__16,linha6_3__15,linha6_3__14,linha6_3__13,linha6_3__12,
              linha6_3__11,linha6_3__10,linha6_3__9,linha6_3__8,linha6_3__7,
              linha6_3__6,linha6_3__5,linha6_3__4,linha6_3__3,linha6_3__2,
              linha6_3__1,linha6_3__0}), .a0 ({linha7_3__63,linha7_3__62,
              linha7_3__61,linha7_3__60,linha7_3__59,linha7_3__58,linha7_3__57,
              linha7_3__56,linha7_3__55,linha7_3__54,linha7_3__53,linha7_3__52,
              linha7_3__51,linha7_3__50,linha7_3__49,linha7_3__48,linha7_3__47,
              linha7_3__46,linha7_3__45,linha7_3__44,linha7_3__43,linha7_3__42,
              linha7_3__41,linha7_3__40,linha7_3__39,linha7_3__38,linha7_3__37,
              linha7_3__36,linha7_3__35,linha7_3__34,linha7_3__33,linha7_3__32,
              linha7_3__31,linha7_3__30,linha7_3__29,linha7_3__28,linha7_3__27,
              linha7_3__26,linha7_3__25,linha7_3__24,linha7_3__23,linha7_3__22,
              linha7_3__21,linha7_3__20,linha7_3__19,linha7_3__18,linha7_3__17,
              linha7_3__16,linha7_3__15,linha7_3__14,linha7_3__13,linha7_3__12,
              linha7_3__11,linha7_3__10,linha7_3__9,linha7_3__8,linha7_3__7,
              linha7_3__6,linha7_3__5,linha7_3__4,linha7_3__3,linha7_3__2,
              linha7_3__1,linha7_3__0}), .s (row_3_rowi_bni3_l)) ;
    juntarComparadores_64 row_4_rowp_bni1_Comp (.g (\$dummy [14]), .l (
                          row_4_rowp_bni1_l), .a ({linha1_2__63,linha1_2__62,
                          linha1_2__61,linha1_2__60,linha1_2__59,linha1_2__58,
                          linha1_2__57,linha1_2__56,linha1_2__55,linha1_2__54,
                          linha1_2__53,linha1_2__52,linha1_2__51,linha1_2__50,
                          linha1_2__49,linha1_2__48,linha1_2__47,linha1_2__46,
                          linha1_2__45,linha1_2__44,linha1_2__43,linha1_2__42,
                          linha1_2__41,linha1_2__40,linha1_2__39,linha1_2__38,
                          linha1_2__37,linha1_2__36,linha1_2__35,linha1_2__34,
                          linha1_2__33,linha1_2__32,linha1_2__31,linha1_2__30,
                          linha1_2__29,linha1_2__28,linha1_2__27,linha1_2__26,
                          linha1_2__25,linha1_2__24,linha1_2__23,linha1_2__22,
                          linha1_2__21,linha1_2__20,linha1_2__19,linha1_2__18,
                          linha1_2__17,linha1_2__16,linha1_2__15,linha1_2__14,
                          linha1_2__13,linha1_2__12,linha1_2__11,linha1_2__10,
                          linha1_2__9,linha1_2__8,linha1_2__7,linha1_2__6,
                          linha1_2__5,linha1_2__4,linha1_2__3,linha1_2__2,
                          linha1_2__1,linha1_2__0}), .b ({linha2_4__63,
                          linha2_4__62,linha2_4__61,linha2_4__60,linha2_4__59,
                          linha2_4__58,linha2_4__57,linha2_4__56,linha2_4__55,
                          linha2_4__54,linha2_4__53,linha2_4__52,linha2_4__51,
                          linha2_4__50,linha2_4__49,linha2_4__48,linha2_4__47,
                          linha2_4__46,linha2_4__45,linha2_4__44,linha2_4__43,
                          linha2_4__42,linha2_4__41,linha2_4__40,linha2_4__39,
                          linha2_4__38,linha2_4__37,linha2_4__36,linha2_4__35,
                          linha2_4__34,linha2_4__33,linha2_4__32,linha2_4__31,
                          linha2_4__30,linha2_4__29,linha2_4__28,linha2_4__27,
                          linha2_4__26,linha2_4__25,linha2_4__24,linha2_4__23,
                          linha2_4__22,linha2_4__21,linha2_4__20,linha2_4__19,
                          linha2_4__18,linha2_4__17,linha2_4__16,linha2_4__15,
                          linha2_4__14,linha2_4__13,linha2_4__12,linha2_4__11,
                          linha2_4__10,linha2_4__9,linha2_4__8,linha2_4__7,
                          linha2_4__6,linha2_4__5,linha2_4__4,linha2_4__3,
                          linha2_4__2,linha2_4__1,linha2_4__0})) ;
    Mux2x1_64 row_4_rowp_bni1_muxMax (.r ({linha1_3__63,linha1_3__62,
              linha1_3__61,linha1_3__60,linha1_3__59,linha1_3__58,linha1_3__57,
              linha1_3__56,linha1_3__55,linha1_3__54,linha1_3__53,linha1_3__52,
              linha1_3__51,linha1_3__50,linha1_3__49,linha1_3__48,linha1_3__47,
              linha1_3__46,linha1_3__45,linha1_3__44,linha1_3__43,linha1_3__42,
              linha1_3__41,linha1_3__40,linha1_3__39,linha1_3__38,linha1_3__37,
              linha1_3__36,linha1_3__35,linha1_3__34,linha1_3__33,linha1_3__32,
              linha1_3__31,linha1_3__30,linha1_3__29,linha1_3__28,linha1_3__27,
              linha1_3__26,linha1_3__25,linha1_3__24,linha1_3__23,linha1_3__22,
              linha1_3__21,linha1_3__20,linha1_3__19,linha1_3__18,linha1_3__17,
              linha1_3__16,linha1_3__15,linha1_3__14,linha1_3__13,linha1_3__12,
              linha1_3__11,linha1_3__10,linha1_3__9,linha1_3__8,linha1_3__7,
              linha1_3__6,linha1_3__5,linha1_3__4,linha1_3__3,linha1_3__2,
              linha1_3__1,linha1_3__0}), .a1 ({linha2_4__63,linha2_4__62,
              linha2_4__61,linha2_4__60,linha2_4__59,linha2_4__58,linha2_4__57,
              linha2_4__56,linha2_4__55,linha2_4__54,linha2_4__53,linha2_4__52,
              linha2_4__51,linha2_4__50,linha2_4__49,linha2_4__48,linha2_4__47,
              linha2_4__46,linha2_4__45,linha2_4__44,linha2_4__43,linha2_4__42,
              linha2_4__41,linha2_4__40,linha2_4__39,linha2_4__38,linha2_4__37,
              linha2_4__36,linha2_4__35,linha2_4__34,linha2_4__33,linha2_4__32,
              linha2_4__31,linha2_4__30,linha2_4__29,linha2_4__28,linha2_4__27,
              linha2_4__26,linha2_4__25,linha2_4__24,linha2_4__23,linha2_4__22,
              linha2_4__21,linha2_4__20,linha2_4__19,linha2_4__18,linha2_4__17,
              linha2_4__16,linha2_4__15,linha2_4__14,linha2_4__13,linha2_4__12,
              linha2_4__11,linha2_4__10,linha2_4__9,linha2_4__8,linha2_4__7,
              linha2_4__6,linha2_4__5,linha2_4__4,linha2_4__3,linha2_4__2,
              linha2_4__1,linha2_4__0}), .a0 ({linha1_2__63,linha1_2__62,
              linha1_2__61,linha1_2__60,linha1_2__59,linha1_2__58,linha1_2__57,
              linha1_2__56,linha1_2__55,linha1_2__54,linha1_2__53,linha1_2__52,
              linha1_2__51,linha1_2__50,linha1_2__49,linha1_2__48,linha1_2__47,
              linha1_2__46,linha1_2__45,linha1_2__44,linha1_2__43,linha1_2__42,
              linha1_2__41,linha1_2__40,linha1_2__39,linha1_2__38,linha1_2__37,
              linha1_2__36,linha1_2__35,linha1_2__34,linha1_2__33,linha1_2__32,
              linha1_2__31,linha1_2__30,linha1_2__29,linha1_2__28,linha1_2__27,
              linha1_2__26,linha1_2__25,linha1_2__24,linha1_2__23,linha1_2__22,
              linha1_2__21,linha1_2__20,linha1_2__19,linha1_2__18,linha1_2__17,
              linha1_2__16,linha1_2__15,linha1_2__14,linha1_2__13,linha1_2__12,
              linha1_2__11,linha1_2__10,linha1_2__9,linha1_2__8,linha1_2__7,
              linha1_2__6,linha1_2__5,linha1_2__4,linha1_2__3,linha1_2__2,
              linha1_2__1,linha1_2__0}), .s (row_4_rowp_bni1_l)) ;
    Mux2x1_64 row_4_rowp_bni1_muxMin (.r ({linha2_5__63,linha2_5__62,
              linha2_5__61,linha2_5__60,linha2_5__59,linha2_5__58,linha2_5__57,
              linha2_5__56,linha2_5__55,linha2_5__54,linha2_5__53,linha2_5__52,
              linha2_5__51,linha2_5__50,linha2_5__49,linha2_5__48,linha2_5__47,
              linha2_5__46,linha2_5__45,linha2_5__44,linha2_5__43,linha2_5__42,
              linha2_5__41,linha2_5__40,linha2_5__39,linha2_5__38,linha2_5__37,
              linha2_5__36,linha2_5__35,linha2_5__34,linha2_5__33,linha2_5__32,
              linha2_5__31,linha2_5__30,linha2_5__29,linha2_5__28,linha2_5__27,
              linha2_5__26,linha2_5__25,linha2_5__24,linha2_5__23,linha2_5__22,
              linha2_5__21,linha2_5__20,linha2_5__19,linha2_5__18,linha2_5__17,
              linha2_5__16,linha2_5__15,linha2_5__14,linha2_5__13,linha2_5__12,
              linha2_5__11,linha2_5__10,linha2_5__9,linha2_5__8,linha2_5__7,
              linha2_5__6,linha2_5__5,linha2_5__4,linha2_5__3,linha2_5__2,
              linha2_5__1,linha2_5__0}), .a1 ({linha1_2__63,linha1_2__62,
              linha1_2__61,linha1_2__60,linha1_2__59,linha1_2__58,linha1_2__57,
              linha1_2__56,linha1_2__55,linha1_2__54,linha1_2__53,linha1_2__52,
              linha1_2__51,linha1_2__50,linha1_2__49,linha1_2__48,linha1_2__47,
              linha1_2__46,linha1_2__45,linha1_2__44,linha1_2__43,linha1_2__42,
              linha1_2__41,linha1_2__40,linha1_2__39,linha1_2__38,linha1_2__37,
              linha1_2__36,linha1_2__35,linha1_2__34,linha1_2__33,linha1_2__32,
              linha1_2__31,linha1_2__30,linha1_2__29,linha1_2__28,linha1_2__27,
              linha1_2__26,linha1_2__25,linha1_2__24,linha1_2__23,linha1_2__22,
              linha1_2__21,linha1_2__20,linha1_2__19,linha1_2__18,linha1_2__17,
              linha1_2__16,linha1_2__15,linha1_2__14,linha1_2__13,linha1_2__12,
              linha1_2__11,linha1_2__10,linha1_2__9,linha1_2__8,linha1_2__7,
              linha1_2__6,linha1_2__5,linha1_2__4,linha1_2__3,linha1_2__2,
              linha1_2__1,linha1_2__0}), .a0 ({linha2_4__63,linha2_4__62,
              linha2_4__61,linha2_4__60,linha2_4__59,linha2_4__58,linha2_4__57,
              linha2_4__56,linha2_4__55,linha2_4__54,linha2_4__53,linha2_4__52,
              linha2_4__51,linha2_4__50,linha2_4__49,linha2_4__48,linha2_4__47,
              linha2_4__46,linha2_4__45,linha2_4__44,linha2_4__43,linha2_4__42,
              linha2_4__41,linha2_4__40,linha2_4__39,linha2_4__38,linha2_4__37,
              linha2_4__36,linha2_4__35,linha2_4__34,linha2_4__33,linha2_4__32,
              linha2_4__31,linha2_4__30,linha2_4__29,linha2_4__28,linha2_4__27,
              linha2_4__26,linha2_4__25,linha2_4__24,linha2_4__23,linha2_4__22,
              linha2_4__21,linha2_4__20,linha2_4__19,linha2_4__18,linha2_4__17,
              linha2_4__16,linha2_4__15,linha2_4__14,linha2_4__13,linha2_4__12,
              linha2_4__11,linha2_4__10,linha2_4__9,linha2_4__8,linha2_4__7,
              linha2_4__6,linha2_4__5,linha2_4__4,linha2_4__3,linha2_4__2,
              linha2_4__1,linha2_4__0}), .s (row_4_rowp_bni1_l)) ;
    juntarComparadores_64 row_4_rowp_bni2_Comp (.g (\$dummy [15]), .l (
                          row_4_rowp_bni2_l), .a ({linha3_4__63,linha3_4__62,
                          linha3_4__61,linha3_4__60,linha3_4__59,linha3_4__58,
                          linha3_4__57,linha3_4__56,linha3_4__55,linha3_4__54,
                          linha3_4__53,linha3_4__52,linha3_4__51,linha3_4__50,
                          linha3_4__49,linha3_4__48,linha3_4__47,linha3_4__46,
                          linha3_4__45,linha3_4__44,linha3_4__43,linha3_4__42,
                          linha3_4__41,linha3_4__40,linha3_4__39,linha3_4__38,
                          linha3_4__37,linha3_4__36,linha3_4__35,linha3_4__34,
                          linha3_4__33,linha3_4__32,linha3_4__31,linha3_4__30,
                          linha3_4__29,linha3_4__28,linha3_4__27,linha3_4__26,
                          linha3_4__25,linha3_4__24,linha3_4__23,linha3_4__22,
                          linha3_4__21,linha3_4__20,linha3_4__19,linha3_4__18,
                          linha3_4__17,linha3_4__16,linha3_4__15,linha3_4__14,
                          linha3_4__13,linha3_4__12,linha3_4__11,linha3_4__10,
                          linha3_4__9,linha3_4__8,linha3_4__7,linha3_4__6,
                          linha3_4__5,linha3_4__4,linha3_4__3,linha3_4__2,
                          linha3_4__1,linha3_4__0}), .b ({linha4_4__63,
                          linha4_4__62,linha4_4__61,linha4_4__60,linha4_4__59,
                          linha4_4__58,linha4_4__57,linha4_4__56,linha4_4__55,
                          linha4_4__54,linha4_4__53,linha4_4__52,linha4_4__51,
                          linha4_4__50,linha4_4__49,linha4_4__48,linha4_4__47,
                          linha4_4__46,linha4_4__45,linha4_4__44,linha4_4__43,
                          linha4_4__42,linha4_4__41,linha4_4__40,linha4_4__39,
                          linha4_4__38,linha4_4__37,linha4_4__36,linha4_4__35,
                          linha4_4__34,linha4_4__33,linha4_4__32,linha4_4__31,
                          linha4_4__30,linha4_4__29,linha4_4__28,linha4_4__27,
                          linha4_4__26,linha4_4__25,linha4_4__24,linha4_4__23,
                          linha4_4__22,linha4_4__21,linha4_4__20,linha4_4__19,
                          linha4_4__18,linha4_4__17,linha4_4__16,linha4_4__15,
                          linha4_4__14,linha4_4__13,linha4_4__12,linha4_4__11,
                          linha4_4__10,linha4_4__9,linha4_4__8,linha4_4__7,
                          linha4_4__6,linha4_4__5,linha4_4__4,linha4_4__3,
                          linha4_4__2,linha4_4__1,linha4_4__0})) ;
    Mux2x1_64 row_4_rowp_bni2_muxMax (.r ({linha3_5__63,linha3_5__62,
              linha3_5__61,linha3_5__60,linha3_5__59,linha3_5__58,linha3_5__57,
              linha3_5__56,linha3_5__55,linha3_5__54,linha3_5__53,linha3_5__52,
              linha3_5__51,linha3_5__50,linha3_5__49,linha3_5__48,linha3_5__47,
              linha3_5__46,linha3_5__45,linha3_5__44,linha3_5__43,linha3_5__42,
              linha3_5__41,linha3_5__40,linha3_5__39,linha3_5__38,linha3_5__37,
              linha3_5__36,linha3_5__35,linha3_5__34,linha3_5__33,linha3_5__32,
              linha3_5__31,linha3_5__30,linha3_5__29,linha3_5__28,linha3_5__27,
              linha3_5__26,linha3_5__25,linha3_5__24,linha3_5__23,linha3_5__22,
              linha3_5__21,linha3_5__20,linha3_5__19,linha3_5__18,linha3_5__17,
              linha3_5__16,linha3_5__15,linha3_5__14,linha3_5__13,linha3_5__12,
              linha3_5__11,linha3_5__10,linha3_5__9,linha3_5__8,linha3_5__7,
              linha3_5__6,linha3_5__5,linha3_5__4,linha3_5__3,linha3_5__2,
              linha3_5__1,linha3_5__0}), .a1 ({linha4_4__63,linha4_4__62,
              linha4_4__61,linha4_4__60,linha4_4__59,linha4_4__58,linha4_4__57,
              linha4_4__56,linha4_4__55,linha4_4__54,linha4_4__53,linha4_4__52,
              linha4_4__51,linha4_4__50,linha4_4__49,linha4_4__48,linha4_4__47,
              linha4_4__46,linha4_4__45,linha4_4__44,linha4_4__43,linha4_4__42,
              linha4_4__41,linha4_4__40,linha4_4__39,linha4_4__38,linha4_4__37,
              linha4_4__36,linha4_4__35,linha4_4__34,linha4_4__33,linha4_4__32,
              linha4_4__31,linha4_4__30,linha4_4__29,linha4_4__28,linha4_4__27,
              linha4_4__26,linha4_4__25,linha4_4__24,linha4_4__23,linha4_4__22,
              linha4_4__21,linha4_4__20,linha4_4__19,linha4_4__18,linha4_4__17,
              linha4_4__16,linha4_4__15,linha4_4__14,linha4_4__13,linha4_4__12,
              linha4_4__11,linha4_4__10,linha4_4__9,linha4_4__8,linha4_4__7,
              linha4_4__6,linha4_4__5,linha4_4__4,linha4_4__3,linha4_4__2,
              linha4_4__1,linha4_4__0}), .a0 ({linha3_4__63,linha3_4__62,
              linha3_4__61,linha3_4__60,linha3_4__59,linha3_4__58,linha3_4__57,
              linha3_4__56,linha3_4__55,linha3_4__54,linha3_4__53,linha3_4__52,
              linha3_4__51,linha3_4__50,linha3_4__49,linha3_4__48,linha3_4__47,
              linha3_4__46,linha3_4__45,linha3_4__44,linha3_4__43,linha3_4__42,
              linha3_4__41,linha3_4__40,linha3_4__39,linha3_4__38,linha3_4__37,
              linha3_4__36,linha3_4__35,linha3_4__34,linha3_4__33,linha3_4__32,
              linha3_4__31,linha3_4__30,linha3_4__29,linha3_4__28,linha3_4__27,
              linha3_4__26,linha3_4__25,linha3_4__24,linha3_4__23,linha3_4__22,
              linha3_4__21,linha3_4__20,linha3_4__19,linha3_4__18,linha3_4__17,
              linha3_4__16,linha3_4__15,linha3_4__14,linha3_4__13,linha3_4__12,
              linha3_4__11,linha3_4__10,linha3_4__9,linha3_4__8,linha3_4__7,
              linha3_4__6,linha3_4__5,linha3_4__4,linha3_4__3,linha3_4__2,
              linha3_4__1,linha3_4__0}), .s (row_4_rowp_bni2_l)) ;
    Mux2x1_64 row_4_rowp_bni2_muxMin (.r ({linha4_5__63,linha4_5__62,
              linha4_5__61,linha4_5__60,linha4_5__59,linha4_5__58,linha4_5__57,
              linha4_5__56,linha4_5__55,linha4_5__54,linha4_5__53,linha4_5__52,
              linha4_5__51,linha4_5__50,linha4_5__49,linha4_5__48,linha4_5__47,
              linha4_5__46,linha4_5__45,linha4_5__44,linha4_5__43,linha4_5__42,
              linha4_5__41,linha4_5__40,linha4_5__39,linha4_5__38,linha4_5__37,
              linha4_5__36,linha4_5__35,linha4_5__34,linha4_5__33,linha4_5__32,
              linha4_5__31,linha4_5__30,linha4_5__29,linha4_5__28,linha4_5__27,
              linha4_5__26,linha4_5__25,linha4_5__24,linha4_5__23,linha4_5__22,
              linha4_5__21,linha4_5__20,linha4_5__19,linha4_5__18,linha4_5__17,
              linha4_5__16,linha4_5__15,linha4_5__14,linha4_5__13,linha4_5__12,
              linha4_5__11,linha4_5__10,linha4_5__9,linha4_5__8,linha4_5__7,
              linha4_5__6,linha4_5__5,linha4_5__4,linha4_5__3,linha4_5__2,
              linha4_5__1,linha4_5__0}), .a1 ({linha3_4__63,linha3_4__62,
              linha3_4__61,linha3_4__60,linha3_4__59,linha3_4__58,linha3_4__57,
              linha3_4__56,linha3_4__55,linha3_4__54,linha3_4__53,linha3_4__52,
              linha3_4__51,linha3_4__50,linha3_4__49,linha3_4__48,linha3_4__47,
              linha3_4__46,linha3_4__45,linha3_4__44,linha3_4__43,linha3_4__42,
              linha3_4__41,linha3_4__40,linha3_4__39,linha3_4__38,linha3_4__37,
              linha3_4__36,linha3_4__35,linha3_4__34,linha3_4__33,linha3_4__32,
              linha3_4__31,linha3_4__30,linha3_4__29,linha3_4__28,linha3_4__27,
              linha3_4__26,linha3_4__25,linha3_4__24,linha3_4__23,linha3_4__22,
              linha3_4__21,linha3_4__20,linha3_4__19,linha3_4__18,linha3_4__17,
              linha3_4__16,linha3_4__15,linha3_4__14,linha3_4__13,linha3_4__12,
              linha3_4__11,linha3_4__10,linha3_4__9,linha3_4__8,linha3_4__7,
              linha3_4__6,linha3_4__5,linha3_4__4,linha3_4__3,linha3_4__2,
              linha3_4__1,linha3_4__0}), .a0 ({linha4_4__63,linha4_4__62,
              linha4_4__61,linha4_4__60,linha4_4__59,linha4_4__58,linha4_4__57,
              linha4_4__56,linha4_4__55,linha4_4__54,linha4_4__53,linha4_4__52,
              linha4_4__51,linha4_4__50,linha4_4__49,linha4_4__48,linha4_4__47,
              linha4_4__46,linha4_4__45,linha4_4__44,linha4_4__43,linha4_4__42,
              linha4_4__41,linha4_4__40,linha4_4__39,linha4_4__38,linha4_4__37,
              linha4_4__36,linha4_4__35,linha4_4__34,linha4_4__33,linha4_4__32,
              linha4_4__31,linha4_4__30,linha4_4__29,linha4_4__28,linha4_4__27,
              linha4_4__26,linha4_4__25,linha4_4__24,linha4_4__23,linha4_4__22,
              linha4_4__21,linha4_4__20,linha4_4__19,linha4_4__18,linha4_4__17,
              linha4_4__16,linha4_4__15,linha4_4__14,linha4_4__13,linha4_4__12,
              linha4_4__11,linha4_4__10,linha4_4__9,linha4_4__8,linha4_4__7,
              linha4_4__6,linha4_4__5,linha4_4__4,linha4_4__3,linha4_4__2,
              linha4_4__1,linha4_4__0}), .s (row_4_rowp_bni2_l)) ;
    juntarComparadores_64 row_4_rowp_bni3_Comp (.g (\$dummy [16]), .l (
                          row_4_rowp_bni3_l), .a ({linha5_4__63,linha5_4__62,
                          linha5_4__61,linha5_4__60,linha5_4__59,linha5_4__58,
                          linha5_4__57,linha5_4__56,linha5_4__55,linha5_4__54,
                          linha5_4__53,linha5_4__52,linha5_4__51,linha5_4__50,
                          linha5_4__49,linha5_4__48,linha5_4__47,linha5_4__46,
                          linha5_4__45,linha5_4__44,linha5_4__43,linha5_4__42,
                          linha5_4__41,linha5_4__40,linha5_4__39,linha5_4__38,
                          linha5_4__37,linha5_4__36,linha5_4__35,linha5_4__34,
                          linha5_4__33,linha5_4__32,linha5_4__31,linha5_4__30,
                          linha5_4__29,linha5_4__28,linha5_4__27,linha5_4__26,
                          linha5_4__25,linha5_4__24,linha5_4__23,linha5_4__22,
                          linha5_4__21,linha5_4__20,linha5_4__19,linha5_4__18,
                          linha5_4__17,linha5_4__16,linha5_4__15,linha5_4__14,
                          linha5_4__13,linha5_4__12,linha5_4__11,linha5_4__10,
                          linha5_4__9,linha5_4__8,linha5_4__7,linha5_4__6,
                          linha5_4__5,linha5_4__4,linha5_4__3,linha5_4__2,
                          linha5_4__1,linha5_4__0}), .b ({linha6_4__63,
                          linha6_4__62,linha6_4__61,linha6_4__60,linha6_4__59,
                          linha6_4__58,linha6_4__57,linha6_4__56,linha6_4__55,
                          linha6_4__54,linha6_4__53,linha6_4__52,linha6_4__51,
                          linha6_4__50,linha6_4__49,linha6_4__48,linha6_4__47,
                          linha6_4__46,linha6_4__45,linha6_4__44,linha6_4__43,
                          linha6_4__42,linha6_4__41,linha6_4__40,linha6_4__39,
                          linha6_4__38,linha6_4__37,linha6_4__36,linha6_4__35,
                          linha6_4__34,linha6_4__33,linha6_4__32,linha6_4__31,
                          linha6_4__30,linha6_4__29,linha6_4__28,linha6_4__27,
                          linha6_4__26,linha6_4__25,linha6_4__24,linha6_4__23,
                          linha6_4__22,linha6_4__21,linha6_4__20,linha6_4__19,
                          linha6_4__18,linha6_4__17,linha6_4__16,linha6_4__15,
                          linha6_4__14,linha6_4__13,linha6_4__12,linha6_4__11,
                          linha6_4__10,linha6_4__9,linha6_4__8,linha6_4__7,
                          linha6_4__6,linha6_4__5,linha6_4__4,linha6_4__3,
                          linha6_4__2,linha6_4__1,linha6_4__0})) ;
    Mux2x1_64 row_4_rowp_bni3_muxMax (.r ({linha5_5__63,linha5_5__62,
              linha5_5__61,linha5_5__60,linha5_5__59,linha5_5__58,linha5_5__57,
              linha5_5__56,linha5_5__55,linha5_5__54,linha5_5__53,linha5_5__52,
              linha5_5__51,linha5_5__50,linha5_5__49,linha5_5__48,linha5_5__47,
              linha5_5__46,linha5_5__45,linha5_5__44,linha5_5__43,linha5_5__42,
              linha5_5__41,linha5_5__40,linha5_5__39,linha5_5__38,linha5_5__37,
              linha5_5__36,linha5_5__35,linha5_5__34,linha5_5__33,linha5_5__32,
              linha5_5__31,linha5_5__30,linha5_5__29,linha5_5__28,linha5_5__27,
              linha5_5__26,linha5_5__25,linha5_5__24,linha5_5__23,linha5_5__22,
              linha5_5__21,linha5_5__20,linha5_5__19,linha5_5__18,linha5_5__17,
              linha5_5__16,linha5_5__15,linha5_5__14,linha5_5__13,linha5_5__12,
              linha5_5__11,linha5_5__10,linha5_5__9,linha5_5__8,linha5_5__7,
              linha5_5__6,linha5_5__5,linha5_5__4,linha5_5__3,linha5_5__2,
              linha5_5__1,linha5_5__0}), .a1 ({linha6_4__63,linha6_4__62,
              linha6_4__61,linha6_4__60,linha6_4__59,linha6_4__58,linha6_4__57,
              linha6_4__56,linha6_4__55,linha6_4__54,linha6_4__53,linha6_4__52,
              linha6_4__51,linha6_4__50,linha6_4__49,linha6_4__48,linha6_4__47,
              linha6_4__46,linha6_4__45,linha6_4__44,linha6_4__43,linha6_4__42,
              linha6_4__41,linha6_4__40,linha6_4__39,linha6_4__38,linha6_4__37,
              linha6_4__36,linha6_4__35,linha6_4__34,linha6_4__33,linha6_4__32,
              linha6_4__31,linha6_4__30,linha6_4__29,linha6_4__28,linha6_4__27,
              linha6_4__26,linha6_4__25,linha6_4__24,linha6_4__23,linha6_4__22,
              linha6_4__21,linha6_4__20,linha6_4__19,linha6_4__18,linha6_4__17,
              linha6_4__16,linha6_4__15,linha6_4__14,linha6_4__13,linha6_4__12,
              linha6_4__11,linha6_4__10,linha6_4__9,linha6_4__8,linha6_4__7,
              linha6_4__6,linha6_4__5,linha6_4__4,linha6_4__3,linha6_4__2,
              linha6_4__1,linha6_4__0}), .a0 ({linha5_4__63,linha5_4__62,
              linha5_4__61,linha5_4__60,linha5_4__59,linha5_4__58,linha5_4__57,
              linha5_4__56,linha5_4__55,linha5_4__54,linha5_4__53,linha5_4__52,
              linha5_4__51,linha5_4__50,linha5_4__49,linha5_4__48,linha5_4__47,
              linha5_4__46,linha5_4__45,linha5_4__44,linha5_4__43,linha5_4__42,
              linha5_4__41,linha5_4__40,linha5_4__39,linha5_4__38,linha5_4__37,
              linha5_4__36,linha5_4__35,linha5_4__34,linha5_4__33,linha5_4__32,
              linha5_4__31,linha5_4__30,linha5_4__29,linha5_4__28,linha5_4__27,
              linha5_4__26,linha5_4__25,linha5_4__24,linha5_4__23,linha5_4__22,
              linha5_4__21,linha5_4__20,linha5_4__19,linha5_4__18,linha5_4__17,
              linha5_4__16,linha5_4__15,linha5_4__14,linha5_4__13,linha5_4__12,
              linha5_4__11,linha5_4__10,linha5_4__9,linha5_4__8,linha5_4__7,
              linha5_4__6,linha5_4__5,linha5_4__4,linha5_4__3,linha5_4__2,
              linha5_4__1,linha5_4__0}), .s (row_4_rowp_bni3_l)) ;
    Mux2x1_64 row_4_rowp_bni3_muxMin (.r ({linha6_5__63,linha6_5__62,
              linha6_5__61,linha6_5__60,linha6_5__59,linha6_5__58,linha6_5__57,
              linha6_5__56,linha6_5__55,linha6_5__54,linha6_5__53,linha6_5__52,
              linha6_5__51,linha6_5__50,linha6_5__49,linha6_5__48,linha6_5__47,
              linha6_5__46,linha6_5__45,linha6_5__44,linha6_5__43,linha6_5__42,
              linha6_5__41,linha6_5__40,linha6_5__39,linha6_5__38,linha6_5__37,
              linha6_5__36,linha6_5__35,linha6_5__34,linha6_5__33,linha6_5__32,
              linha6_5__31,linha6_5__30,linha6_5__29,linha6_5__28,linha6_5__27,
              linha6_5__26,linha6_5__25,linha6_5__24,linha6_5__23,linha6_5__22,
              linha6_5__21,linha6_5__20,linha6_5__19,linha6_5__18,linha6_5__17,
              linha6_5__16,linha6_5__15,linha6_5__14,linha6_5__13,linha6_5__12,
              linha6_5__11,linha6_5__10,linha6_5__9,linha6_5__8,linha6_5__7,
              linha6_5__6,linha6_5__5,linha6_5__4,linha6_5__3,linha6_5__2,
              linha6_5__1,linha6_5__0}), .a1 ({linha5_4__63,linha5_4__62,
              linha5_4__61,linha5_4__60,linha5_4__59,linha5_4__58,linha5_4__57,
              linha5_4__56,linha5_4__55,linha5_4__54,linha5_4__53,linha5_4__52,
              linha5_4__51,linha5_4__50,linha5_4__49,linha5_4__48,linha5_4__47,
              linha5_4__46,linha5_4__45,linha5_4__44,linha5_4__43,linha5_4__42,
              linha5_4__41,linha5_4__40,linha5_4__39,linha5_4__38,linha5_4__37,
              linha5_4__36,linha5_4__35,linha5_4__34,linha5_4__33,linha5_4__32,
              linha5_4__31,linha5_4__30,linha5_4__29,linha5_4__28,linha5_4__27,
              linha5_4__26,linha5_4__25,linha5_4__24,linha5_4__23,linha5_4__22,
              linha5_4__21,linha5_4__20,linha5_4__19,linha5_4__18,linha5_4__17,
              linha5_4__16,linha5_4__15,linha5_4__14,linha5_4__13,linha5_4__12,
              linha5_4__11,linha5_4__10,linha5_4__9,linha5_4__8,linha5_4__7,
              linha5_4__6,linha5_4__5,linha5_4__4,linha5_4__3,linha5_4__2,
              linha5_4__1,linha5_4__0}), .a0 ({linha6_4__63,linha6_4__62,
              linha6_4__61,linha6_4__60,linha6_4__59,linha6_4__58,linha6_4__57,
              linha6_4__56,linha6_4__55,linha6_4__54,linha6_4__53,linha6_4__52,
              linha6_4__51,linha6_4__50,linha6_4__49,linha6_4__48,linha6_4__47,
              linha6_4__46,linha6_4__45,linha6_4__44,linha6_4__43,linha6_4__42,
              linha6_4__41,linha6_4__40,linha6_4__39,linha6_4__38,linha6_4__37,
              linha6_4__36,linha6_4__35,linha6_4__34,linha6_4__33,linha6_4__32,
              linha6_4__31,linha6_4__30,linha6_4__29,linha6_4__28,linha6_4__27,
              linha6_4__26,linha6_4__25,linha6_4__24,linha6_4__23,linha6_4__22,
              linha6_4__21,linha6_4__20,linha6_4__19,linha6_4__18,linha6_4__17,
              linha6_4__16,linha6_4__15,linha6_4__14,linha6_4__13,linha6_4__12,
              linha6_4__11,linha6_4__10,linha6_4__9,linha6_4__8,linha6_4__7,
              linha6_4__6,linha6_4__5,linha6_4__4,linha6_4__3,linha6_4__2,
              linha6_4__1,linha6_4__0}), .s (row_4_rowp_bni3_l)) ;
    juntarComparadores_64 row_4_rowp_bni4_Comp (.g (\$dummy [17]), .l (
                          row_4_rowp_bni4_l), .a ({linha7_4__63,linha7_4__62,
                          linha7_4__61,linha7_4__60,linha7_4__59,linha7_4__58,
                          linha7_4__57,linha7_4__56,linha7_4__55,linha7_4__54,
                          linha7_4__53,linha7_4__52,linha7_4__51,linha7_4__50,
                          linha7_4__49,linha7_4__48,linha7_4__47,linha7_4__46,
                          linha7_4__45,linha7_4__44,linha7_4__43,linha7_4__42,
                          linha7_4__41,linha7_4__40,linha7_4__39,linha7_4__38,
                          linha7_4__37,linha7_4__36,linha7_4__35,linha7_4__34,
                          linha7_4__33,linha7_4__32,linha7_4__31,linha7_4__30,
                          linha7_4__29,linha7_4__28,linha7_4__27,linha7_4__26,
                          linha7_4__25,linha7_4__24,linha7_4__23,linha7_4__22,
                          linha7_4__21,linha7_4__20,linha7_4__19,linha7_4__18,
                          linha7_4__17,linha7_4__16,linha7_4__15,linha7_4__14,
                          linha7_4__13,linha7_4__12,linha7_4__11,linha7_4__10,
                          linha7_4__9,linha7_4__8,linha7_4__7,linha7_4__6,
                          linha7_4__5,linha7_4__4,linha7_4__3,linha7_4__2,
                          linha7_4__1,linha7_4__0}), .b ({linha8_2__63,
                          linha8_2__62,linha8_2__61,linha8_2__60,linha8_2__59,
                          linha8_2__58,linha8_2__57,linha8_2__56,linha8_2__55,
                          linha8_2__54,linha8_2__53,linha8_2__52,linha8_2__51,
                          linha8_2__50,linha8_2__49,linha8_2__48,linha8_2__47,
                          linha8_2__46,linha8_2__45,linha8_2__44,linha8_2__43,
                          linha8_2__42,linha8_2__41,linha8_2__40,linha8_2__39,
                          linha8_2__38,linha8_2__37,linha8_2__36,linha8_2__35,
                          linha8_2__34,linha8_2__33,linha8_2__32,linha8_2__31,
                          linha8_2__30,linha8_2__29,linha8_2__28,linha8_2__27,
                          linha8_2__26,linha8_2__25,linha8_2__24,linha8_2__23,
                          linha8_2__22,linha8_2__21,linha8_2__20,linha8_2__19,
                          linha8_2__18,linha8_2__17,linha8_2__16,linha8_2__15,
                          linha8_2__14,linha8_2__13,linha8_2__12,linha8_2__11,
                          linha8_2__10,linha8_2__9,linha8_2__8,linha8_2__7,
                          linha8_2__6,linha8_2__5,linha8_2__4,linha8_2__3,
                          linha8_2__2,linha8_2__1,linha8_2__0})) ;
    Mux2x1_64 row_4_rowp_bni4_muxMax (.r ({linha7_5__63,linha7_5__62,
              linha7_5__61,linha7_5__60,linha7_5__59,linha7_5__58,linha7_5__57,
              linha7_5__56,linha7_5__55,linha7_5__54,linha7_5__53,linha7_5__52,
              linha7_5__51,linha7_5__50,linha7_5__49,linha7_5__48,linha7_5__47,
              linha7_5__46,linha7_5__45,linha7_5__44,linha7_5__43,linha7_5__42,
              linha7_5__41,linha7_5__40,linha7_5__39,linha7_5__38,linha7_5__37,
              linha7_5__36,linha7_5__35,linha7_5__34,linha7_5__33,linha7_5__32,
              linha7_5__31,linha7_5__30,linha7_5__29,linha7_5__28,linha7_5__27,
              linha7_5__26,linha7_5__25,linha7_5__24,linha7_5__23,linha7_5__22,
              linha7_5__21,linha7_5__20,linha7_5__19,linha7_5__18,linha7_5__17,
              linha7_5__16,linha7_5__15,linha7_5__14,linha7_5__13,linha7_5__12,
              linha7_5__11,linha7_5__10,linha7_5__9,linha7_5__8,linha7_5__7,
              linha7_5__6,linha7_5__5,linha7_5__4,linha7_5__3,linha7_5__2,
              linha7_5__1,linha7_5__0}), .a1 ({linha8_2__63,linha8_2__62,
              linha8_2__61,linha8_2__60,linha8_2__59,linha8_2__58,linha8_2__57,
              linha8_2__56,linha8_2__55,linha8_2__54,linha8_2__53,linha8_2__52,
              linha8_2__51,linha8_2__50,linha8_2__49,linha8_2__48,linha8_2__47,
              linha8_2__46,linha8_2__45,linha8_2__44,linha8_2__43,linha8_2__42,
              linha8_2__41,linha8_2__40,linha8_2__39,linha8_2__38,linha8_2__37,
              linha8_2__36,linha8_2__35,linha8_2__34,linha8_2__33,linha8_2__32,
              linha8_2__31,linha8_2__30,linha8_2__29,linha8_2__28,linha8_2__27,
              linha8_2__26,linha8_2__25,linha8_2__24,linha8_2__23,linha8_2__22,
              linha8_2__21,linha8_2__20,linha8_2__19,linha8_2__18,linha8_2__17,
              linha8_2__16,linha8_2__15,linha8_2__14,linha8_2__13,linha8_2__12,
              linha8_2__11,linha8_2__10,linha8_2__9,linha8_2__8,linha8_2__7,
              linha8_2__6,linha8_2__5,linha8_2__4,linha8_2__3,linha8_2__2,
              linha8_2__1,linha8_2__0}), .a0 ({linha7_4__63,linha7_4__62,
              linha7_4__61,linha7_4__60,linha7_4__59,linha7_4__58,linha7_4__57,
              linha7_4__56,linha7_4__55,linha7_4__54,linha7_4__53,linha7_4__52,
              linha7_4__51,linha7_4__50,linha7_4__49,linha7_4__48,linha7_4__47,
              linha7_4__46,linha7_4__45,linha7_4__44,linha7_4__43,linha7_4__42,
              linha7_4__41,linha7_4__40,linha7_4__39,linha7_4__38,linha7_4__37,
              linha7_4__36,linha7_4__35,linha7_4__34,linha7_4__33,linha7_4__32,
              linha7_4__31,linha7_4__30,linha7_4__29,linha7_4__28,linha7_4__27,
              linha7_4__26,linha7_4__25,linha7_4__24,linha7_4__23,linha7_4__22,
              linha7_4__21,linha7_4__20,linha7_4__19,linha7_4__18,linha7_4__17,
              linha7_4__16,linha7_4__15,linha7_4__14,linha7_4__13,linha7_4__12,
              linha7_4__11,linha7_4__10,linha7_4__9,linha7_4__8,linha7_4__7,
              linha7_4__6,linha7_4__5,linha7_4__4,linha7_4__3,linha7_4__2,
              linha7_4__1,linha7_4__0}), .s (row_4_rowp_bni4_l)) ;
    Mux2x1_64 row_4_rowp_bni4_muxMin (.r ({linha8_3__63,linha8_3__62,
              linha8_3__61,linha8_3__60,linha8_3__59,linha8_3__58,linha8_3__57,
              linha8_3__56,linha8_3__55,linha8_3__54,linha8_3__53,linha8_3__52,
              linha8_3__51,linha8_3__50,linha8_3__49,linha8_3__48,linha8_3__47,
              linha8_3__46,linha8_3__45,linha8_3__44,linha8_3__43,linha8_3__42,
              linha8_3__41,linha8_3__40,linha8_3__39,linha8_3__38,linha8_3__37,
              linha8_3__36,linha8_3__35,linha8_3__34,linha8_3__33,linha8_3__32,
              linha8_3__31,linha8_3__30,linha8_3__29,linha8_3__28,linha8_3__27,
              linha8_3__26,linha8_3__25,linha8_3__24,linha8_3__23,linha8_3__22,
              linha8_3__21,linha8_3__20,linha8_3__19,linha8_3__18,linha8_3__17,
              linha8_3__16,linha8_3__15,linha8_3__14,linha8_3__13,linha8_3__12,
              linha8_3__11,linha8_3__10,linha8_3__9,linha8_3__8,linha8_3__7,
              linha8_3__6,linha8_3__5,linha8_3__4,linha8_3__3,linha8_3__2,
              linha8_3__1,linha8_3__0}), .a1 ({linha7_4__63,linha7_4__62,
              linha7_4__61,linha7_4__60,linha7_4__59,linha7_4__58,linha7_4__57,
              linha7_4__56,linha7_4__55,linha7_4__54,linha7_4__53,linha7_4__52,
              linha7_4__51,linha7_4__50,linha7_4__49,linha7_4__48,linha7_4__47,
              linha7_4__46,linha7_4__45,linha7_4__44,linha7_4__43,linha7_4__42,
              linha7_4__41,linha7_4__40,linha7_4__39,linha7_4__38,linha7_4__37,
              linha7_4__36,linha7_4__35,linha7_4__34,linha7_4__33,linha7_4__32,
              linha7_4__31,linha7_4__30,linha7_4__29,linha7_4__28,linha7_4__27,
              linha7_4__26,linha7_4__25,linha7_4__24,linha7_4__23,linha7_4__22,
              linha7_4__21,linha7_4__20,linha7_4__19,linha7_4__18,linha7_4__17,
              linha7_4__16,linha7_4__15,linha7_4__14,linha7_4__13,linha7_4__12,
              linha7_4__11,linha7_4__10,linha7_4__9,linha7_4__8,linha7_4__7,
              linha7_4__6,linha7_4__5,linha7_4__4,linha7_4__3,linha7_4__2,
              linha7_4__1,linha7_4__0}), .a0 ({linha8_2__63,linha8_2__62,
              linha8_2__61,linha8_2__60,linha8_2__59,linha8_2__58,linha8_2__57,
              linha8_2__56,linha8_2__55,linha8_2__54,linha8_2__53,linha8_2__52,
              linha8_2__51,linha8_2__50,linha8_2__49,linha8_2__48,linha8_2__47,
              linha8_2__46,linha8_2__45,linha8_2__44,linha8_2__43,linha8_2__42,
              linha8_2__41,linha8_2__40,linha8_2__39,linha8_2__38,linha8_2__37,
              linha8_2__36,linha8_2__35,linha8_2__34,linha8_2__33,linha8_2__32,
              linha8_2__31,linha8_2__30,linha8_2__29,linha8_2__28,linha8_2__27,
              linha8_2__26,linha8_2__25,linha8_2__24,linha8_2__23,linha8_2__22,
              linha8_2__21,linha8_2__20,linha8_2__19,linha8_2__18,linha8_2__17,
              linha8_2__16,linha8_2__15,linha8_2__14,linha8_2__13,linha8_2__12,
              linha8_2__11,linha8_2__10,linha8_2__9,linha8_2__8,linha8_2__7,
              linha8_2__6,linha8_2__5,linha8_2__4,linha8_2__3,linha8_2__2,
              linha8_2__1,linha8_2__0}), .s (row_4_rowp_bni4_l)) ;
    juntarComparadores_64 row_5_rowi_bni1_Comp (.g (\$dummy [18]), .l (
                          row_5_rowi_bni1_l), .a ({linha2_5__63,linha2_5__62,
                          linha2_5__61,linha2_5__60,linha2_5__59,linha2_5__58,
                          linha2_5__57,linha2_5__56,linha2_5__55,linha2_5__54,
                          linha2_5__53,linha2_5__52,linha2_5__51,linha2_5__50,
                          linha2_5__49,linha2_5__48,linha2_5__47,linha2_5__46,
                          linha2_5__45,linha2_5__44,linha2_5__43,linha2_5__42,
                          linha2_5__41,linha2_5__40,linha2_5__39,linha2_5__38,
                          linha2_5__37,linha2_5__36,linha2_5__35,linha2_5__34,
                          linha2_5__33,linha2_5__32,linha2_5__31,linha2_5__30,
                          linha2_5__29,linha2_5__28,linha2_5__27,linha2_5__26,
                          linha2_5__25,linha2_5__24,linha2_5__23,linha2_5__22,
                          linha2_5__21,linha2_5__20,linha2_5__19,linha2_5__18,
                          linha2_5__17,linha2_5__16,linha2_5__15,linha2_5__14,
                          linha2_5__13,linha2_5__12,linha2_5__11,linha2_5__10,
                          linha2_5__9,linha2_5__8,linha2_5__7,linha2_5__6,
                          linha2_5__5,linha2_5__4,linha2_5__3,linha2_5__2,
                          linha2_5__1,linha2_5__0}), .b ({linha3_5__63,
                          linha3_5__62,linha3_5__61,linha3_5__60,linha3_5__59,
                          linha3_5__58,linha3_5__57,linha3_5__56,linha3_5__55,
                          linha3_5__54,linha3_5__53,linha3_5__52,linha3_5__51,
                          linha3_5__50,linha3_5__49,linha3_5__48,linha3_5__47,
                          linha3_5__46,linha3_5__45,linha3_5__44,linha3_5__43,
                          linha3_5__42,linha3_5__41,linha3_5__40,linha3_5__39,
                          linha3_5__38,linha3_5__37,linha3_5__36,linha3_5__35,
                          linha3_5__34,linha3_5__33,linha3_5__32,linha3_5__31,
                          linha3_5__30,linha3_5__29,linha3_5__28,linha3_5__27,
                          linha3_5__26,linha3_5__25,linha3_5__24,linha3_5__23,
                          linha3_5__22,linha3_5__21,linha3_5__20,linha3_5__19,
                          linha3_5__18,linha3_5__17,linha3_5__16,linha3_5__15,
                          linha3_5__14,linha3_5__13,linha3_5__12,linha3_5__11,
                          linha3_5__10,linha3_5__9,linha3_5__8,linha3_5__7,
                          linha3_5__6,linha3_5__5,linha3_5__4,linha3_5__3,
                          linha3_5__2,linha3_5__1,linha3_5__0})) ;
    Mux2x1_64 row_5_rowi_bni1_muxMax (.r ({linha2_6__63,linha2_6__62,
              linha2_6__61,linha2_6__60,linha2_6__59,linha2_6__58,linha2_6__57,
              linha2_6__56,linha2_6__55,linha2_6__54,linha2_6__53,linha2_6__52,
              linha2_6__51,linha2_6__50,linha2_6__49,linha2_6__48,linha2_6__47,
              linha2_6__46,linha2_6__45,linha2_6__44,linha2_6__43,linha2_6__42,
              linha2_6__41,linha2_6__40,linha2_6__39,linha2_6__38,linha2_6__37,
              linha2_6__36,linha2_6__35,linha2_6__34,linha2_6__33,linha2_6__32,
              linha2_6__31,linha2_6__30,linha2_6__29,linha2_6__28,linha2_6__27,
              linha2_6__26,linha2_6__25,linha2_6__24,linha2_6__23,linha2_6__22,
              linha2_6__21,linha2_6__20,linha2_6__19,linha2_6__18,linha2_6__17,
              linha2_6__16,linha2_6__15,linha2_6__14,linha2_6__13,linha2_6__12,
              linha2_6__11,linha2_6__10,linha2_6__9,linha2_6__8,linha2_6__7,
              linha2_6__6,linha2_6__5,linha2_6__4,linha2_6__3,linha2_6__2,
              linha2_6__1,linha2_6__0}), .a1 ({linha3_5__63,linha3_5__62,
              linha3_5__61,linha3_5__60,linha3_5__59,linha3_5__58,linha3_5__57,
              linha3_5__56,linha3_5__55,linha3_5__54,linha3_5__53,linha3_5__52,
              linha3_5__51,linha3_5__50,linha3_5__49,linha3_5__48,linha3_5__47,
              linha3_5__46,linha3_5__45,linha3_5__44,linha3_5__43,linha3_5__42,
              linha3_5__41,linha3_5__40,linha3_5__39,linha3_5__38,linha3_5__37,
              linha3_5__36,linha3_5__35,linha3_5__34,linha3_5__33,linha3_5__32,
              linha3_5__31,linha3_5__30,linha3_5__29,linha3_5__28,linha3_5__27,
              linha3_5__26,linha3_5__25,linha3_5__24,linha3_5__23,linha3_5__22,
              linha3_5__21,linha3_5__20,linha3_5__19,linha3_5__18,linha3_5__17,
              linha3_5__16,linha3_5__15,linha3_5__14,linha3_5__13,linha3_5__12,
              linha3_5__11,linha3_5__10,linha3_5__9,linha3_5__8,linha3_5__7,
              linha3_5__6,linha3_5__5,linha3_5__4,linha3_5__3,linha3_5__2,
              linha3_5__1,linha3_5__0}), .a0 ({linha2_5__63,linha2_5__62,
              linha2_5__61,linha2_5__60,linha2_5__59,linha2_5__58,linha2_5__57,
              linha2_5__56,linha2_5__55,linha2_5__54,linha2_5__53,linha2_5__52,
              linha2_5__51,linha2_5__50,linha2_5__49,linha2_5__48,linha2_5__47,
              linha2_5__46,linha2_5__45,linha2_5__44,linha2_5__43,linha2_5__42,
              linha2_5__41,linha2_5__40,linha2_5__39,linha2_5__38,linha2_5__37,
              linha2_5__36,linha2_5__35,linha2_5__34,linha2_5__33,linha2_5__32,
              linha2_5__31,linha2_5__30,linha2_5__29,linha2_5__28,linha2_5__27,
              linha2_5__26,linha2_5__25,linha2_5__24,linha2_5__23,linha2_5__22,
              linha2_5__21,linha2_5__20,linha2_5__19,linha2_5__18,linha2_5__17,
              linha2_5__16,linha2_5__15,linha2_5__14,linha2_5__13,linha2_5__12,
              linha2_5__11,linha2_5__10,linha2_5__9,linha2_5__8,linha2_5__7,
              linha2_5__6,linha2_5__5,linha2_5__4,linha2_5__3,linha2_5__2,
              linha2_5__1,linha2_5__0}), .s (row_5_rowi_bni1_l)) ;
    Mux2x1_64 row_5_rowi_bni1_muxMin (.r ({linha3_6__63,linha3_6__62,
              linha3_6__61,linha3_6__60,linha3_6__59,linha3_6__58,linha3_6__57,
              linha3_6__56,linha3_6__55,linha3_6__54,linha3_6__53,linha3_6__52,
              linha3_6__51,linha3_6__50,linha3_6__49,linha3_6__48,linha3_6__47,
              linha3_6__46,linha3_6__45,linha3_6__44,linha3_6__43,linha3_6__42,
              linha3_6__41,linha3_6__40,linha3_6__39,linha3_6__38,linha3_6__37,
              linha3_6__36,linha3_6__35,linha3_6__34,linha3_6__33,linha3_6__32,
              linha3_6__31,linha3_6__30,linha3_6__29,linha3_6__28,linha3_6__27,
              linha3_6__26,linha3_6__25,linha3_6__24,linha3_6__23,linha3_6__22,
              linha3_6__21,linha3_6__20,linha3_6__19,linha3_6__18,linha3_6__17,
              linha3_6__16,linha3_6__15,linha3_6__14,linha3_6__13,linha3_6__12,
              linha3_6__11,linha3_6__10,linha3_6__9,linha3_6__8,linha3_6__7,
              linha3_6__6,linha3_6__5,linha3_6__4,linha3_6__3,linha3_6__2,
              linha3_6__1,linha3_6__0}), .a1 ({linha2_5__63,linha2_5__62,
              linha2_5__61,linha2_5__60,linha2_5__59,linha2_5__58,linha2_5__57,
              linha2_5__56,linha2_5__55,linha2_5__54,linha2_5__53,linha2_5__52,
              linha2_5__51,linha2_5__50,linha2_5__49,linha2_5__48,linha2_5__47,
              linha2_5__46,linha2_5__45,linha2_5__44,linha2_5__43,linha2_5__42,
              linha2_5__41,linha2_5__40,linha2_5__39,linha2_5__38,linha2_5__37,
              linha2_5__36,linha2_5__35,linha2_5__34,linha2_5__33,linha2_5__32,
              linha2_5__31,linha2_5__30,linha2_5__29,linha2_5__28,linha2_5__27,
              linha2_5__26,linha2_5__25,linha2_5__24,linha2_5__23,linha2_5__22,
              linha2_5__21,linha2_5__20,linha2_5__19,linha2_5__18,linha2_5__17,
              linha2_5__16,linha2_5__15,linha2_5__14,linha2_5__13,linha2_5__12,
              linha2_5__11,linha2_5__10,linha2_5__9,linha2_5__8,linha2_5__7,
              linha2_5__6,linha2_5__5,linha2_5__4,linha2_5__3,linha2_5__2,
              linha2_5__1,linha2_5__0}), .a0 ({linha3_5__63,linha3_5__62,
              linha3_5__61,linha3_5__60,linha3_5__59,linha3_5__58,linha3_5__57,
              linha3_5__56,linha3_5__55,linha3_5__54,linha3_5__53,linha3_5__52,
              linha3_5__51,linha3_5__50,linha3_5__49,linha3_5__48,linha3_5__47,
              linha3_5__46,linha3_5__45,linha3_5__44,linha3_5__43,linha3_5__42,
              linha3_5__41,linha3_5__40,linha3_5__39,linha3_5__38,linha3_5__37,
              linha3_5__36,linha3_5__35,linha3_5__34,linha3_5__33,linha3_5__32,
              linha3_5__31,linha3_5__30,linha3_5__29,linha3_5__28,linha3_5__27,
              linha3_5__26,linha3_5__25,linha3_5__24,linha3_5__23,linha3_5__22,
              linha3_5__21,linha3_5__20,linha3_5__19,linha3_5__18,linha3_5__17,
              linha3_5__16,linha3_5__15,linha3_5__14,linha3_5__13,linha3_5__12,
              linha3_5__11,linha3_5__10,linha3_5__9,linha3_5__8,linha3_5__7,
              linha3_5__6,linha3_5__5,linha3_5__4,linha3_5__3,linha3_5__2,
              linha3_5__1,linha3_5__0}), .s (row_5_rowi_bni1_l)) ;
    juntarComparadores_64 row_5_rowi_bni2_Comp (.g (\$dummy [19]), .l (
                          row_5_rowi_bni2_l), .a ({linha4_5__63,linha4_5__62,
                          linha4_5__61,linha4_5__60,linha4_5__59,linha4_5__58,
                          linha4_5__57,linha4_5__56,linha4_5__55,linha4_5__54,
                          linha4_5__53,linha4_5__52,linha4_5__51,linha4_5__50,
                          linha4_5__49,linha4_5__48,linha4_5__47,linha4_5__46,
                          linha4_5__45,linha4_5__44,linha4_5__43,linha4_5__42,
                          linha4_5__41,linha4_5__40,linha4_5__39,linha4_5__38,
                          linha4_5__37,linha4_5__36,linha4_5__35,linha4_5__34,
                          linha4_5__33,linha4_5__32,linha4_5__31,linha4_5__30,
                          linha4_5__29,linha4_5__28,linha4_5__27,linha4_5__26,
                          linha4_5__25,linha4_5__24,linha4_5__23,linha4_5__22,
                          linha4_5__21,linha4_5__20,linha4_5__19,linha4_5__18,
                          linha4_5__17,linha4_5__16,linha4_5__15,linha4_5__14,
                          linha4_5__13,linha4_5__12,linha4_5__11,linha4_5__10,
                          linha4_5__9,linha4_5__8,linha4_5__7,linha4_5__6,
                          linha4_5__5,linha4_5__4,linha4_5__3,linha4_5__2,
                          linha4_5__1,linha4_5__0}), .b ({linha5_5__63,
                          linha5_5__62,linha5_5__61,linha5_5__60,linha5_5__59,
                          linha5_5__58,linha5_5__57,linha5_5__56,linha5_5__55,
                          linha5_5__54,linha5_5__53,linha5_5__52,linha5_5__51,
                          linha5_5__50,linha5_5__49,linha5_5__48,linha5_5__47,
                          linha5_5__46,linha5_5__45,linha5_5__44,linha5_5__43,
                          linha5_5__42,linha5_5__41,linha5_5__40,linha5_5__39,
                          linha5_5__38,linha5_5__37,linha5_5__36,linha5_5__35,
                          linha5_5__34,linha5_5__33,linha5_5__32,linha5_5__31,
                          linha5_5__30,linha5_5__29,linha5_5__28,linha5_5__27,
                          linha5_5__26,linha5_5__25,linha5_5__24,linha5_5__23,
                          linha5_5__22,linha5_5__21,linha5_5__20,linha5_5__19,
                          linha5_5__18,linha5_5__17,linha5_5__16,linha5_5__15,
                          linha5_5__14,linha5_5__13,linha5_5__12,linha5_5__11,
                          linha5_5__10,linha5_5__9,linha5_5__8,linha5_5__7,
                          linha5_5__6,linha5_5__5,linha5_5__4,linha5_5__3,
                          linha5_5__2,linha5_5__1,linha5_5__0})) ;
    Mux2x1_64 row_5_rowi_bni2_muxMax (.r ({linha4_6__63,linha4_6__62,
              linha4_6__61,linha4_6__60,linha4_6__59,linha4_6__58,linha4_6__57,
              linha4_6__56,linha4_6__55,linha4_6__54,linha4_6__53,linha4_6__52,
              linha4_6__51,linha4_6__50,linha4_6__49,linha4_6__48,linha4_6__47,
              linha4_6__46,linha4_6__45,linha4_6__44,linha4_6__43,linha4_6__42,
              linha4_6__41,linha4_6__40,linha4_6__39,linha4_6__38,linha4_6__37,
              linha4_6__36,linha4_6__35,linha4_6__34,linha4_6__33,linha4_6__32,
              linha4_6__31,linha4_6__30,linha4_6__29,linha4_6__28,linha4_6__27,
              linha4_6__26,linha4_6__25,linha4_6__24,linha4_6__23,linha4_6__22,
              linha4_6__21,linha4_6__20,linha4_6__19,linha4_6__18,linha4_6__17,
              linha4_6__16,linha4_6__15,linha4_6__14,linha4_6__13,linha4_6__12,
              linha4_6__11,linha4_6__10,linha4_6__9,linha4_6__8,linha4_6__7,
              linha4_6__6,linha4_6__5,linha4_6__4,linha4_6__3,linha4_6__2,
              linha4_6__1,linha4_6__0}), .a1 ({linha5_5__63,linha5_5__62,
              linha5_5__61,linha5_5__60,linha5_5__59,linha5_5__58,linha5_5__57,
              linha5_5__56,linha5_5__55,linha5_5__54,linha5_5__53,linha5_5__52,
              linha5_5__51,linha5_5__50,linha5_5__49,linha5_5__48,linha5_5__47,
              linha5_5__46,linha5_5__45,linha5_5__44,linha5_5__43,linha5_5__42,
              linha5_5__41,linha5_5__40,linha5_5__39,linha5_5__38,linha5_5__37,
              linha5_5__36,linha5_5__35,linha5_5__34,linha5_5__33,linha5_5__32,
              linha5_5__31,linha5_5__30,linha5_5__29,linha5_5__28,linha5_5__27,
              linha5_5__26,linha5_5__25,linha5_5__24,linha5_5__23,linha5_5__22,
              linha5_5__21,linha5_5__20,linha5_5__19,linha5_5__18,linha5_5__17,
              linha5_5__16,linha5_5__15,linha5_5__14,linha5_5__13,linha5_5__12,
              linha5_5__11,linha5_5__10,linha5_5__9,linha5_5__8,linha5_5__7,
              linha5_5__6,linha5_5__5,linha5_5__4,linha5_5__3,linha5_5__2,
              linha5_5__1,linha5_5__0}), .a0 ({linha4_5__63,linha4_5__62,
              linha4_5__61,linha4_5__60,linha4_5__59,linha4_5__58,linha4_5__57,
              linha4_5__56,linha4_5__55,linha4_5__54,linha4_5__53,linha4_5__52,
              linha4_5__51,linha4_5__50,linha4_5__49,linha4_5__48,linha4_5__47,
              linha4_5__46,linha4_5__45,linha4_5__44,linha4_5__43,linha4_5__42,
              linha4_5__41,linha4_5__40,linha4_5__39,linha4_5__38,linha4_5__37,
              linha4_5__36,linha4_5__35,linha4_5__34,linha4_5__33,linha4_5__32,
              linha4_5__31,linha4_5__30,linha4_5__29,linha4_5__28,linha4_5__27,
              linha4_5__26,linha4_5__25,linha4_5__24,linha4_5__23,linha4_5__22,
              linha4_5__21,linha4_5__20,linha4_5__19,linha4_5__18,linha4_5__17,
              linha4_5__16,linha4_5__15,linha4_5__14,linha4_5__13,linha4_5__12,
              linha4_5__11,linha4_5__10,linha4_5__9,linha4_5__8,linha4_5__7,
              linha4_5__6,linha4_5__5,linha4_5__4,linha4_5__3,linha4_5__2,
              linha4_5__1,linha4_5__0}), .s (row_5_rowi_bni2_l)) ;
    Mux2x1_64 row_5_rowi_bni2_muxMin (.r ({linha5_6__63,linha5_6__62,
              linha5_6__61,linha5_6__60,linha5_6__59,linha5_6__58,linha5_6__57,
              linha5_6__56,linha5_6__55,linha5_6__54,linha5_6__53,linha5_6__52,
              linha5_6__51,linha5_6__50,linha5_6__49,linha5_6__48,linha5_6__47,
              linha5_6__46,linha5_6__45,linha5_6__44,linha5_6__43,linha5_6__42,
              linha5_6__41,linha5_6__40,linha5_6__39,linha5_6__38,linha5_6__37,
              linha5_6__36,linha5_6__35,linha5_6__34,linha5_6__33,linha5_6__32,
              linha5_6__31,linha5_6__30,linha5_6__29,linha5_6__28,linha5_6__27,
              linha5_6__26,linha5_6__25,linha5_6__24,linha5_6__23,linha5_6__22,
              linha5_6__21,linha5_6__20,linha5_6__19,linha5_6__18,linha5_6__17,
              linha5_6__16,linha5_6__15,linha5_6__14,linha5_6__13,linha5_6__12,
              linha5_6__11,linha5_6__10,linha5_6__9,linha5_6__8,linha5_6__7,
              linha5_6__6,linha5_6__5,linha5_6__4,linha5_6__3,linha5_6__2,
              linha5_6__1,linha5_6__0}), .a1 ({linha4_5__63,linha4_5__62,
              linha4_5__61,linha4_5__60,linha4_5__59,linha4_5__58,linha4_5__57,
              linha4_5__56,linha4_5__55,linha4_5__54,linha4_5__53,linha4_5__52,
              linha4_5__51,linha4_5__50,linha4_5__49,linha4_5__48,linha4_5__47,
              linha4_5__46,linha4_5__45,linha4_5__44,linha4_5__43,linha4_5__42,
              linha4_5__41,linha4_5__40,linha4_5__39,linha4_5__38,linha4_5__37,
              linha4_5__36,linha4_5__35,linha4_5__34,linha4_5__33,linha4_5__32,
              linha4_5__31,linha4_5__30,linha4_5__29,linha4_5__28,linha4_5__27,
              linha4_5__26,linha4_5__25,linha4_5__24,linha4_5__23,linha4_5__22,
              linha4_5__21,linha4_5__20,linha4_5__19,linha4_5__18,linha4_5__17,
              linha4_5__16,linha4_5__15,linha4_5__14,linha4_5__13,linha4_5__12,
              linha4_5__11,linha4_5__10,linha4_5__9,linha4_5__8,linha4_5__7,
              linha4_5__6,linha4_5__5,linha4_5__4,linha4_5__3,linha4_5__2,
              linha4_5__1,linha4_5__0}), .a0 ({linha5_5__63,linha5_5__62,
              linha5_5__61,linha5_5__60,linha5_5__59,linha5_5__58,linha5_5__57,
              linha5_5__56,linha5_5__55,linha5_5__54,linha5_5__53,linha5_5__52,
              linha5_5__51,linha5_5__50,linha5_5__49,linha5_5__48,linha5_5__47,
              linha5_5__46,linha5_5__45,linha5_5__44,linha5_5__43,linha5_5__42,
              linha5_5__41,linha5_5__40,linha5_5__39,linha5_5__38,linha5_5__37,
              linha5_5__36,linha5_5__35,linha5_5__34,linha5_5__33,linha5_5__32,
              linha5_5__31,linha5_5__30,linha5_5__29,linha5_5__28,linha5_5__27,
              linha5_5__26,linha5_5__25,linha5_5__24,linha5_5__23,linha5_5__22,
              linha5_5__21,linha5_5__20,linha5_5__19,linha5_5__18,linha5_5__17,
              linha5_5__16,linha5_5__15,linha5_5__14,linha5_5__13,linha5_5__12,
              linha5_5__11,linha5_5__10,linha5_5__9,linha5_5__8,linha5_5__7,
              linha5_5__6,linha5_5__5,linha5_5__4,linha5_5__3,linha5_5__2,
              linha5_5__1,linha5_5__0}), .s (row_5_rowi_bni2_l)) ;
    juntarComparadores_64 row_5_rowi_bni3_Comp (.g (\$dummy [20]), .l (
                          row_5_rowi_bni3_l), .a ({linha6_5__63,linha6_5__62,
                          linha6_5__61,linha6_5__60,linha6_5__59,linha6_5__58,
                          linha6_5__57,linha6_5__56,linha6_5__55,linha6_5__54,
                          linha6_5__53,linha6_5__52,linha6_5__51,linha6_5__50,
                          linha6_5__49,linha6_5__48,linha6_5__47,linha6_5__46,
                          linha6_5__45,linha6_5__44,linha6_5__43,linha6_5__42,
                          linha6_5__41,linha6_5__40,linha6_5__39,linha6_5__38,
                          linha6_5__37,linha6_5__36,linha6_5__35,linha6_5__34,
                          linha6_5__33,linha6_5__32,linha6_5__31,linha6_5__30,
                          linha6_5__29,linha6_5__28,linha6_5__27,linha6_5__26,
                          linha6_5__25,linha6_5__24,linha6_5__23,linha6_5__22,
                          linha6_5__21,linha6_5__20,linha6_5__19,linha6_5__18,
                          linha6_5__17,linha6_5__16,linha6_5__15,linha6_5__14,
                          linha6_5__13,linha6_5__12,linha6_5__11,linha6_5__10,
                          linha6_5__9,linha6_5__8,linha6_5__7,linha6_5__6,
                          linha6_5__5,linha6_5__4,linha6_5__3,linha6_5__2,
                          linha6_5__1,linha6_5__0}), .b ({linha7_5__63,
                          linha7_5__62,linha7_5__61,linha7_5__60,linha7_5__59,
                          linha7_5__58,linha7_5__57,linha7_5__56,linha7_5__55,
                          linha7_5__54,linha7_5__53,linha7_5__52,linha7_5__51,
                          linha7_5__50,linha7_5__49,linha7_5__48,linha7_5__47,
                          linha7_5__46,linha7_5__45,linha7_5__44,linha7_5__43,
                          linha7_5__42,linha7_5__41,linha7_5__40,linha7_5__39,
                          linha7_5__38,linha7_5__37,linha7_5__36,linha7_5__35,
                          linha7_5__34,linha7_5__33,linha7_5__32,linha7_5__31,
                          linha7_5__30,linha7_5__29,linha7_5__28,linha7_5__27,
                          linha7_5__26,linha7_5__25,linha7_5__24,linha7_5__23,
                          linha7_5__22,linha7_5__21,linha7_5__20,linha7_5__19,
                          linha7_5__18,linha7_5__17,linha7_5__16,linha7_5__15,
                          linha7_5__14,linha7_5__13,linha7_5__12,linha7_5__11,
                          linha7_5__10,linha7_5__9,linha7_5__8,linha7_5__7,
                          linha7_5__6,linha7_5__5,linha7_5__4,linha7_5__3,
                          linha7_5__2,linha7_5__1,linha7_5__0})) ;
    Mux2x1_64 row_5_rowi_bni3_muxMax (.r ({linha6_6__63,linha6_6__62,
              linha6_6__61,linha6_6__60,linha6_6__59,linha6_6__58,linha6_6__57,
              linha6_6__56,linha6_6__55,linha6_6__54,linha6_6__53,linha6_6__52,
              linha6_6__51,linha6_6__50,linha6_6__49,linha6_6__48,linha6_6__47,
              linha6_6__46,linha6_6__45,linha6_6__44,linha6_6__43,linha6_6__42,
              linha6_6__41,linha6_6__40,linha6_6__39,linha6_6__38,linha6_6__37,
              linha6_6__36,linha6_6__35,linha6_6__34,linha6_6__33,linha6_6__32,
              linha6_6__31,linha6_6__30,linha6_6__29,linha6_6__28,linha6_6__27,
              linha6_6__26,linha6_6__25,linha6_6__24,linha6_6__23,linha6_6__22,
              linha6_6__21,linha6_6__20,linha6_6__19,linha6_6__18,linha6_6__17,
              linha6_6__16,linha6_6__15,linha6_6__14,linha6_6__13,linha6_6__12,
              linha6_6__11,linha6_6__10,linha6_6__9,linha6_6__8,linha6_6__7,
              linha6_6__6,linha6_6__5,linha6_6__4,linha6_6__3,linha6_6__2,
              linha6_6__1,linha6_6__0}), .a1 ({linha7_5__63,linha7_5__62,
              linha7_5__61,linha7_5__60,linha7_5__59,linha7_5__58,linha7_5__57,
              linha7_5__56,linha7_5__55,linha7_5__54,linha7_5__53,linha7_5__52,
              linha7_5__51,linha7_5__50,linha7_5__49,linha7_5__48,linha7_5__47,
              linha7_5__46,linha7_5__45,linha7_5__44,linha7_5__43,linha7_5__42,
              linha7_5__41,linha7_5__40,linha7_5__39,linha7_5__38,linha7_5__37,
              linha7_5__36,linha7_5__35,linha7_5__34,linha7_5__33,linha7_5__32,
              linha7_5__31,linha7_5__30,linha7_5__29,linha7_5__28,linha7_5__27,
              linha7_5__26,linha7_5__25,linha7_5__24,linha7_5__23,linha7_5__22,
              linha7_5__21,linha7_5__20,linha7_5__19,linha7_5__18,linha7_5__17,
              linha7_5__16,linha7_5__15,linha7_5__14,linha7_5__13,linha7_5__12,
              linha7_5__11,linha7_5__10,linha7_5__9,linha7_5__8,linha7_5__7,
              linha7_5__6,linha7_5__5,linha7_5__4,linha7_5__3,linha7_5__2,
              linha7_5__1,linha7_5__0}), .a0 ({linha6_5__63,linha6_5__62,
              linha6_5__61,linha6_5__60,linha6_5__59,linha6_5__58,linha6_5__57,
              linha6_5__56,linha6_5__55,linha6_5__54,linha6_5__53,linha6_5__52,
              linha6_5__51,linha6_5__50,linha6_5__49,linha6_5__48,linha6_5__47,
              linha6_5__46,linha6_5__45,linha6_5__44,linha6_5__43,linha6_5__42,
              linha6_5__41,linha6_5__40,linha6_5__39,linha6_5__38,linha6_5__37,
              linha6_5__36,linha6_5__35,linha6_5__34,linha6_5__33,linha6_5__32,
              linha6_5__31,linha6_5__30,linha6_5__29,linha6_5__28,linha6_5__27,
              linha6_5__26,linha6_5__25,linha6_5__24,linha6_5__23,linha6_5__22,
              linha6_5__21,linha6_5__20,linha6_5__19,linha6_5__18,linha6_5__17,
              linha6_5__16,linha6_5__15,linha6_5__14,linha6_5__13,linha6_5__12,
              linha6_5__11,linha6_5__10,linha6_5__9,linha6_5__8,linha6_5__7,
              linha6_5__6,linha6_5__5,linha6_5__4,linha6_5__3,linha6_5__2,
              linha6_5__1,linha6_5__0}), .s (row_5_rowi_bni3_l)) ;
    Mux2x1_64 row_5_rowi_bni3_muxMin (.r ({linha7_6__63,linha7_6__62,
              linha7_6__61,linha7_6__60,linha7_6__59,linha7_6__58,linha7_6__57,
              linha7_6__56,linha7_6__55,linha7_6__54,linha7_6__53,linha7_6__52,
              linha7_6__51,linha7_6__50,linha7_6__49,linha7_6__48,linha7_6__47,
              linha7_6__46,linha7_6__45,linha7_6__44,linha7_6__43,linha7_6__42,
              linha7_6__41,linha7_6__40,linha7_6__39,linha7_6__38,linha7_6__37,
              linha7_6__36,linha7_6__35,linha7_6__34,linha7_6__33,linha7_6__32,
              linha7_6__31,linha7_6__30,linha7_6__29,linha7_6__28,linha7_6__27,
              linha7_6__26,linha7_6__25,linha7_6__24,linha7_6__23,linha7_6__22,
              linha7_6__21,linha7_6__20,linha7_6__19,linha7_6__18,linha7_6__17,
              linha7_6__16,linha7_6__15,linha7_6__14,linha7_6__13,linha7_6__12,
              linha7_6__11,linha7_6__10,linha7_6__9,linha7_6__8,linha7_6__7,
              linha7_6__6,linha7_6__5,linha7_6__4,linha7_6__3,linha7_6__2,
              linha7_6__1,linha7_6__0}), .a1 ({linha6_5__63,linha6_5__62,
              linha6_5__61,linha6_5__60,linha6_5__59,linha6_5__58,linha6_5__57,
              linha6_5__56,linha6_5__55,linha6_5__54,linha6_5__53,linha6_5__52,
              linha6_5__51,linha6_5__50,linha6_5__49,linha6_5__48,linha6_5__47,
              linha6_5__46,linha6_5__45,linha6_5__44,linha6_5__43,linha6_5__42,
              linha6_5__41,linha6_5__40,linha6_5__39,linha6_5__38,linha6_5__37,
              linha6_5__36,linha6_5__35,linha6_5__34,linha6_5__33,linha6_5__32,
              linha6_5__31,linha6_5__30,linha6_5__29,linha6_5__28,linha6_5__27,
              linha6_5__26,linha6_5__25,linha6_5__24,linha6_5__23,linha6_5__22,
              linha6_5__21,linha6_5__20,linha6_5__19,linha6_5__18,linha6_5__17,
              linha6_5__16,linha6_5__15,linha6_5__14,linha6_5__13,linha6_5__12,
              linha6_5__11,linha6_5__10,linha6_5__9,linha6_5__8,linha6_5__7,
              linha6_5__6,linha6_5__5,linha6_5__4,linha6_5__3,linha6_5__2,
              linha6_5__1,linha6_5__0}), .a0 ({linha7_5__63,linha7_5__62,
              linha7_5__61,linha7_5__60,linha7_5__59,linha7_5__58,linha7_5__57,
              linha7_5__56,linha7_5__55,linha7_5__54,linha7_5__53,linha7_5__52,
              linha7_5__51,linha7_5__50,linha7_5__49,linha7_5__48,linha7_5__47,
              linha7_5__46,linha7_5__45,linha7_5__44,linha7_5__43,linha7_5__42,
              linha7_5__41,linha7_5__40,linha7_5__39,linha7_5__38,linha7_5__37,
              linha7_5__36,linha7_5__35,linha7_5__34,linha7_5__33,linha7_5__32,
              linha7_5__31,linha7_5__30,linha7_5__29,linha7_5__28,linha7_5__27,
              linha7_5__26,linha7_5__25,linha7_5__24,linha7_5__23,linha7_5__22,
              linha7_5__21,linha7_5__20,linha7_5__19,linha7_5__18,linha7_5__17,
              linha7_5__16,linha7_5__15,linha7_5__14,linha7_5__13,linha7_5__12,
              linha7_5__11,linha7_5__10,linha7_5__9,linha7_5__8,linha7_5__7,
              linha7_5__6,linha7_5__5,linha7_5__4,linha7_5__3,linha7_5__2,
              linha7_5__1,linha7_5__0}), .s (row_5_rowi_bni3_l)) ;
    juntarComparadores_64 row_6_rowp_bni1_Comp (.g (\$dummy [21]), .l (
                          row_6_rowp_bni1_l), .a ({linha1_3__63,linha1_3__62,
                          linha1_3__61,linha1_3__60,linha1_3__59,linha1_3__58,
                          linha1_3__57,linha1_3__56,linha1_3__55,linha1_3__54,
                          linha1_3__53,linha1_3__52,linha1_3__51,linha1_3__50,
                          linha1_3__49,linha1_3__48,linha1_3__47,linha1_3__46,
                          linha1_3__45,linha1_3__44,linha1_3__43,linha1_3__42,
                          linha1_3__41,linha1_3__40,linha1_3__39,linha1_3__38,
                          linha1_3__37,linha1_3__36,linha1_3__35,linha1_3__34,
                          linha1_3__33,linha1_3__32,linha1_3__31,linha1_3__30,
                          linha1_3__29,linha1_3__28,linha1_3__27,linha1_3__26,
                          linha1_3__25,linha1_3__24,linha1_3__23,linha1_3__22,
                          linha1_3__21,linha1_3__20,linha1_3__19,linha1_3__18,
                          linha1_3__17,linha1_3__16,linha1_3__15,linha1_3__14,
                          linha1_3__13,linha1_3__12,linha1_3__11,linha1_3__10,
                          linha1_3__9,linha1_3__8,linha1_3__7,linha1_3__6,
                          linha1_3__5,linha1_3__4,linha1_3__3,linha1_3__2,
                          linha1_3__1,linha1_3__0}), .b ({linha2_6__63,
                          linha2_6__62,linha2_6__61,linha2_6__60,linha2_6__59,
                          linha2_6__58,linha2_6__57,linha2_6__56,linha2_6__55,
                          linha2_6__54,linha2_6__53,linha2_6__52,linha2_6__51,
                          linha2_6__50,linha2_6__49,linha2_6__48,linha2_6__47,
                          linha2_6__46,linha2_6__45,linha2_6__44,linha2_6__43,
                          linha2_6__42,linha2_6__41,linha2_6__40,linha2_6__39,
                          linha2_6__38,linha2_6__37,linha2_6__36,linha2_6__35,
                          linha2_6__34,linha2_6__33,linha2_6__32,linha2_6__31,
                          linha2_6__30,linha2_6__29,linha2_6__28,linha2_6__27,
                          linha2_6__26,linha2_6__25,linha2_6__24,linha2_6__23,
                          linha2_6__22,linha2_6__21,linha2_6__20,linha2_6__19,
                          linha2_6__18,linha2_6__17,linha2_6__16,linha2_6__15,
                          linha2_6__14,linha2_6__13,linha2_6__12,linha2_6__11,
                          linha2_6__10,linha2_6__9,linha2_6__8,linha2_6__7,
                          linha2_6__6,linha2_6__5,linha2_6__4,linha2_6__3,
                          linha2_6__2,linha2_6__1,linha2_6__0})) ;
    Mux2x1_64 row_6_rowp_bni1_muxMax (.r ({y1[63],y1[62],y1[61],y1[60],y1[59],
              y1[58],y1[57],y1[56],y1[55],y1[54],y1[53],y1[52],y1[51],y1[50],
              y1[49],y1[48],y1[47],y1[46],y1[45],y1[44],y1[43],y1[42],y1[41],
              y1[40],y1[39],y1[38],y1[37],y1[36],y1[35],y1[34],y1[33],y1[32],
              y1[31],y1[30],y1[29],y1[28],y1[27],y1[26],y1[25],y1[24],y1[23],
              y1[22],y1[21],y1[20],y1[19],y1[18],y1[17],y1[16],y1[15],y1[14],
              y1[13],y1[12],y1[11],y1[10],y1[9],y1[8],y1[7],y1[6],y1[5],y1[4],
              y1[3],y1[2],y1[1],y1[0]}), .a1 ({linha2_6__63,linha2_6__62,
              linha2_6__61,linha2_6__60,linha2_6__59,linha2_6__58,linha2_6__57,
              linha2_6__56,linha2_6__55,linha2_6__54,linha2_6__53,linha2_6__52,
              linha2_6__51,linha2_6__50,linha2_6__49,linha2_6__48,linha2_6__47,
              linha2_6__46,linha2_6__45,linha2_6__44,linha2_6__43,linha2_6__42,
              linha2_6__41,linha2_6__40,linha2_6__39,linha2_6__38,linha2_6__37,
              linha2_6__36,linha2_6__35,linha2_6__34,linha2_6__33,linha2_6__32,
              linha2_6__31,linha2_6__30,linha2_6__29,linha2_6__28,linha2_6__27,
              linha2_6__26,linha2_6__25,linha2_6__24,linha2_6__23,linha2_6__22,
              linha2_6__21,linha2_6__20,linha2_6__19,linha2_6__18,linha2_6__17,
              linha2_6__16,linha2_6__15,linha2_6__14,linha2_6__13,linha2_6__12,
              linha2_6__11,linha2_6__10,linha2_6__9,linha2_6__8,linha2_6__7,
              linha2_6__6,linha2_6__5,linha2_6__4,linha2_6__3,linha2_6__2,
              linha2_6__1,linha2_6__0}), .a0 ({linha1_3__63,linha1_3__62,
              linha1_3__61,linha1_3__60,linha1_3__59,linha1_3__58,linha1_3__57,
              linha1_3__56,linha1_3__55,linha1_3__54,linha1_3__53,linha1_3__52,
              linha1_3__51,linha1_3__50,linha1_3__49,linha1_3__48,linha1_3__47,
              linha1_3__46,linha1_3__45,linha1_3__44,linha1_3__43,linha1_3__42,
              linha1_3__41,linha1_3__40,linha1_3__39,linha1_3__38,linha1_3__37,
              linha1_3__36,linha1_3__35,linha1_3__34,linha1_3__33,linha1_3__32,
              linha1_3__31,linha1_3__30,linha1_3__29,linha1_3__28,linha1_3__27,
              linha1_3__26,linha1_3__25,linha1_3__24,linha1_3__23,linha1_3__22,
              linha1_3__21,linha1_3__20,linha1_3__19,linha1_3__18,linha1_3__17,
              linha1_3__16,linha1_3__15,linha1_3__14,linha1_3__13,linha1_3__12,
              linha1_3__11,linha1_3__10,linha1_3__9,linha1_3__8,linha1_3__7,
              linha1_3__6,linha1_3__5,linha1_3__4,linha1_3__3,linha1_3__2,
              linha1_3__1,linha1_3__0}), .s (row_6_rowp_bni1_l)) ;
    Mux2x1_64 row_6_rowp_bni1_muxMin (.r ({linha2_7__63,linha2_7__62,
              linha2_7__61,linha2_7__60,linha2_7__59,linha2_7__58,linha2_7__57,
              linha2_7__56,linha2_7__55,linha2_7__54,linha2_7__53,linha2_7__52,
              linha2_7__51,linha2_7__50,linha2_7__49,linha2_7__48,linha2_7__47,
              linha2_7__46,linha2_7__45,linha2_7__44,linha2_7__43,linha2_7__42,
              linha2_7__41,linha2_7__40,linha2_7__39,linha2_7__38,linha2_7__37,
              linha2_7__36,linha2_7__35,linha2_7__34,linha2_7__33,linha2_7__32,
              linha2_7__31,linha2_7__30,linha2_7__29,linha2_7__28,linha2_7__27,
              linha2_7__26,linha2_7__25,linha2_7__24,linha2_7__23,linha2_7__22,
              linha2_7__21,linha2_7__20,linha2_7__19,linha2_7__18,linha2_7__17,
              linha2_7__16,linha2_7__15,linha2_7__14,linha2_7__13,linha2_7__12,
              linha2_7__11,linha2_7__10,linha2_7__9,linha2_7__8,linha2_7__7,
              linha2_7__6,linha2_7__5,linha2_7__4,linha2_7__3,linha2_7__2,
              linha2_7__1,linha2_7__0}), .a1 ({linha1_3__63,linha1_3__62,
              linha1_3__61,linha1_3__60,linha1_3__59,linha1_3__58,linha1_3__57,
              linha1_3__56,linha1_3__55,linha1_3__54,linha1_3__53,linha1_3__52,
              linha1_3__51,linha1_3__50,linha1_3__49,linha1_3__48,linha1_3__47,
              linha1_3__46,linha1_3__45,linha1_3__44,linha1_3__43,linha1_3__42,
              linha1_3__41,linha1_3__40,linha1_3__39,linha1_3__38,linha1_3__37,
              linha1_3__36,linha1_3__35,linha1_3__34,linha1_3__33,linha1_3__32,
              linha1_3__31,linha1_3__30,linha1_3__29,linha1_3__28,linha1_3__27,
              linha1_3__26,linha1_3__25,linha1_3__24,linha1_3__23,linha1_3__22,
              linha1_3__21,linha1_3__20,linha1_3__19,linha1_3__18,linha1_3__17,
              linha1_3__16,linha1_3__15,linha1_3__14,linha1_3__13,linha1_3__12,
              linha1_3__11,linha1_3__10,linha1_3__9,linha1_3__8,linha1_3__7,
              linha1_3__6,linha1_3__5,linha1_3__4,linha1_3__3,linha1_3__2,
              linha1_3__1,linha1_3__0}), .a0 ({linha2_6__63,linha2_6__62,
              linha2_6__61,linha2_6__60,linha2_6__59,linha2_6__58,linha2_6__57,
              linha2_6__56,linha2_6__55,linha2_6__54,linha2_6__53,linha2_6__52,
              linha2_6__51,linha2_6__50,linha2_6__49,linha2_6__48,linha2_6__47,
              linha2_6__46,linha2_6__45,linha2_6__44,linha2_6__43,linha2_6__42,
              linha2_6__41,linha2_6__40,linha2_6__39,linha2_6__38,linha2_6__37,
              linha2_6__36,linha2_6__35,linha2_6__34,linha2_6__33,linha2_6__32,
              linha2_6__31,linha2_6__30,linha2_6__29,linha2_6__28,linha2_6__27,
              linha2_6__26,linha2_6__25,linha2_6__24,linha2_6__23,linha2_6__22,
              linha2_6__21,linha2_6__20,linha2_6__19,linha2_6__18,linha2_6__17,
              linha2_6__16,linha2_6__15,linha2_6__14,linha2_6__13,linha2_6__12,
              linha2_6__11,linha2_6__10,linha2_6__9,linha2_6__8,linha2_6__7,
              linha2_6__6,linha2_6__5,linha2_6__4,linha2_6__3,linha2_6__2,
              linha2_6__1,linha2_6__0}), .s (row_6_rowp_bni1_l)) ;
    juntarComparadores_64 row_6_rowp_bni2_Comp (.g (\$dummy [22]), .l (
                          row_6_rowp_bni2_l), .a ({linha3_6__63,linha3_6__62,
                          linha3_6__61,linha3_6__60,linha3_6__59,linha3_6__58,
                          linha3_6__57,linha3_6__56,linha3_6__55,linha3_6__54,
                          linha3_6__53,linha3_6__52,linha3_6__51,linha3_6__50,
                          linha3_6__49,linha3_6__48,linha3_6__47,linha3_6__46,
                          linha3_6__45,linha3_6__44,linha3_6__43,linha3_6__42,
                          linha3_6__41,linha3_6__40,linha3_6__39,linha3_6__38,
                          linha3_6__37,linha3_6__36,linha3_6__35,linha3_6__34,
                          linha3_6__33,linha3_6__32,linha3_6__31,linha3_6__30,
                          linha3_6__29,linha3_6__28,linha3_6__27,linha3_6__26,
                          linha3_6__25,linha3_6__24,linha3_6__23,linha3_6__22,
                          linha3_6__21,linha3_6__20,linha3_6__19,linha3_6__18,
                          linha3_6__17,linha3_6__16,linha3_6__15,linha3_6__14,
                          linha3_6__13,linha3_6__12,linha3_6__11,linha3_6__10,
                          linha3_6__9,linha3_6__8,linha3_6__7,linha3_6__6,
                          linha3_6__5,linha3_6__4,linha3_6__3,linha3_6__2,
                          linha3_6__1,linha3_6__0}), .b ({linha4_6__63,
                          linha4_6__62,linha4_6__61,linha4_6__60,linha4_6__59,
                          linha4_6__58,linha4_6__57,linha4_6__56,linha4_6__55,
                          linha4_6__54,linha4_6__53,linha4_6__52,linha4_6__51,
                          linha4_6__50,linha4_6__49,linha4_6__48,linha4_6__47,
                          linha4_6__46,linha4_6__45,linha4_6__44,linha4_6__43,
                          linha4_6__42,linha4_6__41,linha4_6__40,linha4_6__39,
                          linha4_6__38,linha4_6__37,linha4_6__36,linha4_6__35,
                          linha4_6__34,linha4_6__33,linha4_6__32,linha4_6__31,
                          linha4_6__30,linha4_6__29,linha4_6__28,linha4_6__27,
                          linha4_6__26,linha4_6__25,linha4_6__24,linha4_6__23,
                          linha4_6__22,linha4_6__21,linha4_6__20,linha4_6__19,
                          linha4_6__18,linha4_6__17,linha4_6__16,linha4_6__15,
                          linha4_6__14,linha4_6__13,linha4_6__12,linha4_6__11,
                          linha4_6__10,linha4_6__9,linha4_6__8,linha4_6__7,
                          linha4_6__6,linha4_6__5,linha4_6__4,linha4_6__3,
                          linha4_6__2,linha4_6__1,linha4_6__0})) ;
    Mux2x1_64 row_6_rowp_bni2_muxMax (.r ({linha3_7__63,linha3_7__62,
              linha3_7__61,linha3_7__60,linha3_7__59,linha3_7__58,linha3_7__57,
              linha3_7__56,linha3_7__55,linha3_7__54,linha3_7__53,linha3_7__52,
              linha3_7__51,linha3_7__50,linha3_7__49,linha3_7__48,linha3_7__47,
              linha3_7__46,linha3_7__45,linha3_7__44,linha3_7__43,linha3_7__42,
              linha3_7__41,linha3_7__40,linha3_7__39,linha3_7__38,linha3_7__37,
              linha3_7__36,linha3_7__35,linha3_7__34,linha3_7__33,linha3_7__32,
              linha3_7__31,linha3_7__30,linha3_7__29,linha3_7__28,linha3_7__27,
              linha3_7__26,linha3_7__25,linha3_7__24,linha3_7__23,linha3_7__22,
              linha3_7__21,linha3_7__20,linha3_7__19,linha3_7__18,linha3_7__17,
              linha3_7__16,linha3_7__15,linha3_7__14,linha3_7__13,linha3_7__12,
              linha3_7__11,linha3_7__10,linha3_7__9,linha3_7__8,linha3_7__7,
              linha3_7__6,linha3_7__5,linha3_7__4,linha3_7__3,linha3_7__2,
              linha3_7__1,linha3_7__0}), .a1 ({linha4_6__63,linha4_6__62,
              linha4_6__61,linha4_6__60,linha4_6__59,linha4_6__58,linha4_6__57,
              linha4_6__56,linha4_6__55,linha4_6__54,linha4_6__53,linha4_6__52,
              linha4_6__51,linha4_6__50,linha4_6__49,linha4_6__48,linha4_6__47,
              linha4_6__46,linha4_6__45,linha4_6__44,linha4_6__43,linha4_6__42,
              linha4_6__41,linha4_6__40,linha4_6__39,linha4_6__38,linha4_6__37,
              linha4_6__36,linha4_6__35,linha4_6__34,linha4_6__33,linha4_6__32,
              linha4_6__31,linha4_6__30,linha4_6__29,linha4_6__28,linha4_6__27,
              linha4_6__26,linha4_6__25,linha4_6__24,linha4_6__23,linha4_6__22,
              linha4_6__21,linha4_6__20,linha4_6__19,linha4_6__18,linha4_6__17,
              linha4_6__16,linha4_6__15,linha4_6__14,linha4_6__13,linha4_6__12,
              linha4_6__11,linha4_6__10,linha4_6__9,linha4_6__8,linha4_6__7,
              linha4_6__6,linha4_6__5,linha4_6__4,linha4_6__3,linha4_6__2,
              linha4_6__1,linha4_6__0}), .a0 ({linha3_6__63,linha3_6__62,
              linha3_6__61,linha3_6__60,linha3_6__59,linha3_6__58,linha3_6__57,
              linha3_6__56,linha3_6__55,linha3_6__54,linha3_6__53,linha3_6__52,
              linha3_6__51,linha3_6__50,linha3_6__49,linha3_6__48,linha3_6__47,
              linha3_6__46,linha3_6__45,linha3_6__44,linha3_6__43,linha3_6__42,
              linha3_6__41,linha3_6__40,linha3_6__39,linha3_6__38,linha3_6__37,
              linha3_6__36,linha3_6__35,linha3_6__34,linha3_6__33,linha3_6__32,
              linha3_6__31,linha3_6__30,linha3_6__29,linha3_6__28,linha3_6__27,
              linha3_6__26,linha3_6__25,linha3_6__24,linha3_6__23,linha3_6__22,
              linha3_6__21,linha3_6__20,linha3_6__19,linha3_6__18,linha3_6__17,
              linha3_6__16,linha3_6__15,linha3_6__14,linha3_6__13,linha3_6__12,
              linha3_6__11,linha3_6__10,linha3_6__9,linha3_6__8,linha3_6__7,
              linha3_6__6,linha3_6__5,linha3_6__4,linha3_6__3,linha3_6__2,
              linha3_6__1,linha3_6__0}), .s (row_6_rowp_bni2_l)) ;
    Mux2x1_64 row_6_rowp_bni2_muxMin (.r ({linha4_7__63,linha4_7__62,
              linha4_7__61,linha4_7__60,linha4_7__59,linha4_7__58,linha4_7__57,
              linha4_7__56,linha4_7__55,linha4_7__54,linha4_7__53,linha4_7__52,
              linha4_7__51,linha4_7__50,linha4_7__49,linha4_7__48,linha4_7__47,
              linha4_7__46,linha4_7__45,linha4_7__44,linha4_7__43,linha4_7__42,
              linha4_7__41,linha4_7__40,linha4_7__39,linha4_7__38,linha4_7__37,
              linha4_7__36,linha4_7__35,linha4_7__34,linha4_7__33,linha4_7__32,
              linha4_7__31,linha4_7__30,linha4_7__29,linha4_7__28,linha4_7__27,
              linha4_7__26,linha4_7__25,linha4_7__24,linha4_7__23,linha4_7__22,
              linha4_7__21,linha4_7__20,linha4_7__19,linha4_7__18,linha4_7__17,
              linha4_7__16,linha4_7__15,linha4_7__14,linha4_7__13,linha4_7__12,
              linha4_7__11,linha4_7__10,linha4_7__9,linha4_7__8,linha4_7__7,
              linha4_7__6,linha4_7__5,linha4_7__4,linha4_7__3,linha4_7__2,
              linha4_7__1,linha4_7__0}), .a1 ({linha3_6__63,linha3_6__62,
              linha3_6__61,linha3_6__60,linha3_6__59,linha3_6__58,linha3_6__57,
              linha3_6__56,linha3_6__55,linha3_6__54,linha3_6__53,linha3_6__52,
              linha3_6__51,linha3_6__50,linha3_6__49,linha3_6__48,linha3_6__47,
              linha3_6__46,linha3_6__45,linha3_6__44,linha3_6__43,linha3_6__42,
              linha3_6__41,linha3_6__40,linha3_6__39,linha3_6__38,linha3_6__37,
              linha3_6__36,linha3_6__35,linha3_6__34,linha3_6__33,linha3_6__32,
              linha3_6__31,linha3_6__30,linha3_6__29,linha3_6__28,linha3_6__27,
              linha3_6__26,linha3_6__25,linha3_6__24,linha3_6__23,linha3_6__22,
              linha3_6__21,linha3_6__20,linha3_6__19,linha3_6__18,linha3_6__17,
              linha3_6__16,linha3_6__15,linha3_6__14,linha3_6__13,linha3_6__12,
              linha3_6__11,linha3_6__10,linha3_6__9,linha3_6__8,linha3_6__7,
              linha3_6__6,linha3_6__5,linha3_6__4,linha3_6__3,linha3_6__2,
              linha3_6__1,linha3_6__0}), .a0 ({linha4_6__63,linha4_6__62,
              linha4_6__61,linha4_6__60,linha4_6__59,linha4_6__58,linha4_6__57,
              linha4_6__56,linha4_6__55,linha4_6__54,linha4_6__53,linha4_6__52,
              linha4_6__51,linha4_6__50,linha4_6__49,linha4_6__48,linha4_6__47,
              linha4_6__46,linha4_6__45,linha4_6__44,linha4_6__43,linha4_6__42,
              linha4_6__41,linha4_6__40,linha4_6__39,linha4_6__38,linha4_6__37,
              linha4_6__36,linha4_6__35,linha4_6__34,linha4_6__33,linha4_6__32,
              linha4_6__31,linha4_6__30,linha4_6__29,linha4_6__28,linha4_6__27,
              linha4_6__26,linha4_6__25,linha4_6__24,linha4_6__23,linha4_6__22,
              linha4_6__21,linha4_6__20,linha4_6__19,linha4_6__18,linha4_6__17,
              linha4_6__16,linha4_6__15,linha4_6__14,linha4_6__13,linha4_6__12,
              linha4_6__11,linha4_6__10,linha4_6__9,linha4_6__8,linha4_6__7,
              linha4_6__6,linha4_6__5,linha4_6__4,linha4_6__3,linha4_6__2,
              linha4_6__1,linha4_6__0}), .s (row_6_rowp_bni2_l)) ;
    juntarComparadores_64 row_6_rowp_bni3_Comp (.g (\$dummy [23]), .l (
                          row_6_rowp_bni3_l), .a ({linha5_6__63,linha5_6__62,
                          linha5_6__61,linha5_6__60,linha5_6__59,linha5_6__58,
                          linha5_6__57,linha5_6__56,linha5_6__55,linha5_6__54,
                          linha5_6__53,linha5_6__52,linha5_6__51,linha5_6__50,
                          linha5_6__49,linha5_6__48,linha5_6__47,linha5_6__46,
                          linha5_6__45,linha5_6__44,linha5_6__43,linha5_6__42,
                          linha5_6__41,linha5_6__40,linha5_6__39,linha5_6__38,
                          linha5_6__37,linha5_6__36,linha5_6__35,linha5_6__34,
                          linha5_6__33,linha5_6__32,linha5_6__31,linha5_6__30,
                          linha5_6__29,linha5_6__28,linha5_6__27,linha5_6__26,
                          linha5_6__25,linha5_6__24,linha5_6__23,linha5_6__22,
                          linha5_6__21,linha5_6__20,linha5_6__19,linha5_6__18,
                          linha5_6__17,linha5_6__16,linha5_6__15,linha5_6__14,
                          linha5_6__13,linha5_6__12,linha5_6__11,linha5_6__10,
                          linha5_6__9,linha5_6__8,linha5_6__7,linha5_6__6,
                          linha5_6__5,linha5_6__4,linha5_6__3,linha5_6__2,
                          linha5_6__1,linha5_6__0}), .b ({linha6_6__63,
                          linha6_6__62,linha6_6__61,linha6_6__60,linha6_6__59,
                          linha6_6__58,linha6_6__57,linha6_6__56,linha6_6__55,
                          linha6_6__54,linha6_6__53,linha6_6__52,linha6_6__51,
                          linha6_6__50,linha6_6__49,linha6_6__48,linha6_6__47,
                          linha6_6__46,linha6_6__45,linha6_6__44,linha6_6__43,
                          linha6_6__42,linha6_6__41,linha6_6__40,linha6_6__39,
                          linha6_6__38,linha6_6__37,linha6_6__36,linha6_6__35,
                          linha6_6__34,linha6_6__33,linha6_6__32,linha6_6__31,
                          linha6_6__30,linha6_6__29,linha6_6__28,linha6_6__27,
                          linha6_6__26,linha6_6__25,linha6_6__24,linha6_6__23,
                          linha6_6__22,linha6_6__21,linha6_6__20,linha6_6__19,
                          linha6_6__18,linha6_6__17,linha6_6__16,linha6_6__15,
                          linha6_6__14,linha6_6__13,linha6_6__12,linha6_6__11,
                          linha6_6__10,linha6_6__9,linha6_6__8,linha6_6__7,
                          linha6_6__6,linha6_6__5,linha6_6__4,linha6_6__3,
                          linha6_6__2,linha6_6__1,linha6_6__0})) ;
    Mux2x1_64 row_6_rowp_bni3_muxMax (.r ({linha5_7__63,linha5_7__62,
              linha5_7__61,linha5_7__60,linha5_7__59,linha5_7__58,linha5_7__57,
              linha5_7__56,linha5_7__55,linha5_7__54,linha5_7__53,linha5_7__52,
              linha5_7__51,linha5_7__50,linha5_7__49,linha5_7__48,linha5_7__47,
              linha5_7__46,linha5_7__45,linha5_7__44,linha5_7__43,linha5_7__42,
              linha5_7__41,linha5_7__40,linha5_7__39,linha5_7__38,linha5_7__37,
              linha5_7__36,linha5_7__35,linha5_7__34,linha5_7__33,linha5_7__32,
              linha5_7__31,linha5_7__30,linha5_7__29,linha5_7__28,linha5_7__27,
              linha5_7__26,linha5_7__25,linha5_7__24,linha5_7__23,linha5_7__22,
              linha5_7__21,linha5_7__20,linha5_7__19,linha5_7__18,linha5_7__17,
              linha5_7__16,linha5_7__15,linha5_7__14,linha5_7__13,linha5_7__12,
              linha5_7__11,linha5_7__10,linha5_7__9,linha5_7__8,linha5_7__7,
              linha5_7__6,linha5_7__5,linha5_7__4,linha5_7__3,linha5_7__2,
              linha5_7__1,linha5_7__0}), .a1 ({linha6_6__63,linha6_6__62,
              linha6_6__61,linha6_6__60,linha6_6__59,linha6_6__58,linha6_6__57,
              linha6_6__56,linha6_6__55,linha6_6__54,linha6_6__53,linha6_6__52,
              linha6_6__51,linha6_6__50,linha6_6__49,linha6_6__48,linha6_6__47,
              linha6_6__46,linha6_6__45,linha6_6__44,linha6_6__43,linha6_6__42,
              linha6_6__41,linha6_6__40,linha6_6__39,linha6_6__38,linha6_6__37,
              linha6_6__36,linha6_6__35,linha6_6__34,linha6_6__33,linha6_6__32,
              linha6_6__31,linha6_6__30,linha6_6__29,linha6_6__28,linha6_6__27,
              linha6_6__26,linha6_6__25,linha6_6__24,linha6_6__23,linha6_6__22,
              linha6_6__21,linha6_6__20,linha6_6__19,linha6_6__18,linha6_6__17,
              linha6_6__16,linha6_6__15,linha6_6__14,linha6_6__13,linha6_6__12,
              linha6_6__11,linha6_6__10,linha6_6__9,linha6_6__8,linha6_6__7,
              linha6_6__6,linha6_6__5,linha6_6__4,linha6_6__3,linha6_6__2,
              linha6_6__1,linha6_6__0}), .a0 ({linha5_6__63,linha5_6__62,
              linha5_6__61,linha5_6__60,linha5_6__59,linha5_6__58,linha5_6__57,
              linha5_6__56,linha5_6__55,linha5_6__54,linha5_6__53,linha5_6__52,
              linha5_6__51,linha5_6__50,linha5_6__49,linha5_6__48,linha5_6__47,
              linha5_6__46,linha5_6__45,linha5_6__44,linha5_6__43,linha5_6__42,
              linha5_6__41,linha5_6__40,linha5_6__39,linha5_6__38,linha5_6__37,
              linha5_6__36,linha5_6__35,linha5_6__34,linha5_6__33,linha5_6__32,
              linha5_6__31,linha5_6__30,linha5_6__29,linha5_6__28,linha5_6__27,
              linha5_6__26,linha5_6__25,linha5_6__24,linha5_6__23,linha5_6__22,
              linha5_6__21,linha5_6__20,linha5_6__19,linha5_6__18,linha5_6__17,
              linha5_6__16,linha5_6__15,linha5_6__14,linha5_6__13,linha5_6__12,
              linha5_6__11,linha5_6__10,linha5_6__9,linha5_6__8,linha5_6__7,
              linha5_6__6,linha5_6__5,linha5_6__4,linha5_6__3,linha5_6__2,
              linha5_6__1,linha5_6__0}), .s (row_6_rowp_bni3_l)) ;
    Mux2x1_64 row_6_rowp_bni3_muxMin (.r ({linha6_7__63,linha6_7__62,
              linha6_7__61,linha6_7__60,linha6_7__59,linha6_7__58,linha6_7__57,
              linha6_7__56,linha6_7__55,linha6_7__54,linha6_7__53,linha6_7__52,
              linha6_7__51,linha6_7__50,linha6_7__49,linha6_7__48,linha6_7__47,
              linha6_7__46,linha6_7__45,linha6_7__44,linha6_7__43,linha6_7__42,
              linha6_7__41,linha6_7__40,linha6_7__39,linha6_7__38,linha6_7__37,
              linha6_7__36,linha6_7__35,linha6_7__34,linha6_7__33,linha6_7__32,
              linha6_7__31,linha6_7__30,linha6_7__29,linha6_7__28,linha6_7__27,
              linha6_7__26,linha6_7__25,linha6_7__24,linha6_7__23,linha6_7__22,
              linha6_7__21,linha6_7__20,linha6_7__19,linha6_7__18,linha6_7__17,
              linha6_7__16,linha6_7__15,linha6_7__14,linha6_7__13,linha6_7__12,
              linha6_7__11,linha6_7__10,linha6_7__9,linha6_7__8,linha6_7__7,
              linha6_7__6,linha6_7__5,linha6_7__4,linha6_7__3,linha6_7__2,
              linha6_7__1,linha6_7__0}), .a1 ({linha5_6__63,linha5_6__62,
              linha5_6__61,linha5_6__60,linha5_6__59,linha5_6__58,linha5_6__57,
              linha5_6__56,linha5_6__55,linha5_6__54,linha5_6__53,linha5_6__52,
              linha5_6__51,linha5_6__50,linha5_6__49,linha5_6__48,linha5_6__47,
              linha5_6__46,linha5_6__45,linha5_6__44,linha5_6__43,linha5_6__42,
              linha5_6__41,linha5_6__40,linha5_6__39,linha5_6__38,linha5_6__37,
              linha5_6__36,linha5_6__35,linha5_6__34,linha5_6__33,linha5_6__32,
              linha5_6__31,linha5_6__30,linha5_6__29,linha5_6__28,linha5_6__27,
              linha5_6__26,linha5_6__25,linha5_6__24,linha5_6__23,linha5_6__22,
              linha5_6__21,linha5_6__20,linha5_6__19,linha5_6__18,linha5_6__17,
              linha5_6__16,linha5_6__15,linha5_6__14,linha5_6__13,linha5_6__12,
              linha5_6__11,linha5_6__10,linha5_6__9,linha5_6__8,linha5_6__7,
              linha5_6__6,linha5_6__5,linha5_6__4,linha5_6__3,linha5_6__2,
              linha5_6__1,linha5_6__0}), .a0 ({linha6_6__63,linha6_6__62,
              linha6_6__61,linha6_6__60,linha6_6__59,linha6_6__58,linha6_6__57,
              linha6_6__56,linha6_6__55,linha6_6__54,linha6_6__53,linha6_6__52,
              linha6_6__51,linha6_6__50,linha6_6__49,linha6_6__48,linha6_6__47,
              linha6_6__46,linha6_6__45,linha6_6__44,linha6_6__43,linha6_6__42,
              linha6_6__41,linha6_6__40,linha6_6__39,linha6_6__38,linha6_6__37,
              linha6_6__36,linha6_6__35,linha6_6__34,linha6_6__33,linha6_6__32,
              linha6_6__31,linha6_6__30,linha6_6__29,linha6_6__28,linha6_6__27,
              linha6_6__26,linha6_6__25,linha6_6__24,linha6_6__23,linha6_6__22,
              linha6_6__21,linha6_6__20,linha6_6__19,linha6_6__18,linha6_6__17,
              linha6_6__16,linha6_6__15,linha6_6__14,linha6_6__13,linha6_6__12,
              linha6_6__11,linha6_6__10,linha6_6__9,linha6_6__8,linha6_6__7,
              linha6_6__6,linha6_6__5,linha6_6__4,linha6_6__3,linha6_6__2,
              linha6_6__1,linha6_6__0}), .s (row_6_rowp_bni3_l)) ;
    juntarComparadores_64 row_6_rowp_bni4_Comp (.g (\$dummy [24]), .l (
                          row_6_rowp_bni4_l), .a ({linha7_6__63,linha7_6__62,
                          linha7_6__61,linha7_6__60,linha7_6__59,linha7_6__58,
                          linha7_6__57,linha7_6__56,linha7_6__55,linha7_6__54,
                          linha7_6__53,linha7_6__52,linha7_6__51,linha7_6__50,
                          linha7_6__49,linha7_6__48,linha7_6__47,linha7_6__46,
                          linha7_6__45,linha7_6__44,linha7_6__43,linha7_6__42,
                          linha7_6__41,linha7_6__40,linha7_6__39,linha7_6__38,
                          linha7_6__37,linha7_6__36,linha7_6__35,linha7_6__34,
                          linha7_6__33,linha7_6__32,linha7_6__31,linha7_6__30,
                          linha7_6__29,linha7_6__28,linha7_6__27,linha7_6__26,
                          linha7_6__25,linha7_6__24,linha7_6__23,linha7_6__22,
                          linha7_6__21,linha7_6__20,linha7_6__19,linha7_6__18,
                          linha7_6__17,linha7_6__16,linha7_6__15,linha7_6__14,
                          linha7_6__13,linha7_6__12,linha7_6__11,linha7_6__10,
                          linha7_6__9,linha7_6__8,linha7_6__7,linha7_6__6,
                          linha7_6__5,linha7_6__4,linha7_6__3,linha7_6__2,
                          linha7_6__1,linha7_6__0}), .b ({linha8_3__63,
                          linha8_3__62,linha8_3__61,linha8_3__60,linha8_3__59,
                          linha8_3__58,linha8_3__57,linha8_3__56,linha8_3__55,
                          linha8_3__54,linha8_3__53,linha8_3__52,linha8_3__51,
                          linha8_3__50,linha8_3__49,linha8_3__48,linha8_3__47,
                          linha8_3__46,linha8_3__45,linha8_3__44,linha8_3__43,
                          linha8_3__42,linha8_3__41,linha8_3__40,linha8_3__39,
                          linha8_3__38,linha8_3__37,linha8_3__36,linha8_3__35,
                          linha8_3__34,linha8_3__33,linha8_3__32,linha8_3__31,
                          linha8_3__30,linha8_3__29,linha8_3__28,linha8_3__27,
                          linha8_3__26,linha8_3__25,linha8_3__24,linha8_3__23,
                          linha8_3__22,linha8_3__21,linha8_3__20,linha8_3__19,
                          linha8_3__18,linha8_3__17,linha8_3__16,linha8_3__15,
                          linha8_3__14,linha8_3__13,linha8_3__12,linha8_3__11,
                          linha8_3__10,linha8_3__9,linha8_3__8,linha8_3__7,
                          linha8_3__6,linha8_3__5,linha8_3__4,linha8_3__3,
                          linha8_3__2,linha8_3__1,linha8_3__0})) ;
    Mux2x1_64 row_6_rowp_bni4_muxMax (.r ({linha7_7__63,linha7_7__62,
              linha7_7__61,linha7_7__60,linha7_7__59,linha7_7__58,linha7_7__57,
              linha7_7__56,linha7_7__55,linha7_7__54,linha7_7__53,linha7_7__52,
              linha7_7__51,linha7_7__50,linha7_7__49,linha7_7__48,linha7_7__47,
              linha7_7__46,linha7_7__45,linha7_7__44,linha7_7__43,linha7_7__42,
              linha7_7__41,linha7_7__40,linha7_7__39,linha7_7__38,linha7_7__37,
              linha7_7__36,linha7_7__35,linha7_7__34,linha7_7__33,linha7_7__32,
              linha7_7__31,linha7_7__30,linha7_7__29,linha7_7__28,linha7_7__27,
              linha7_7__26,linha7_7__25,linha7_7__24,linha7_7__23,linha7_7__22,
              linha7_7__21,linha7_7__20,linha7_7__19,linha7_7__18,linha7_7__17,
              linha7_7__16,linha7_7__15,linha7_7__14,linha7_7__13,linha7_7__12,
              linha7_7__11,linha7_7__10,linha7_7__9,linha7_7__8,linha7_7__7,
              linha7_7__6,linha7_7__5,linha7_7__4,linha7_7__3,linha7_7__2,
              linha7_7__1,linha7_7__0}), .a1 ({linha8_3__63,linha8_3__62,
              linha8_3__61,linha8_3__60,linha8_3__59,linha8_3__58,linha8_3__57,
              linha8_3__56,linha8_3__55,linha8_3__54,linha8_3__53,linha8_3__52,
              linha8_3__51,linha8_3__50,linha8_3__49,linha8_3__48,linha8_3__47,
              linha8_3__46,linha8_3__45,linha8_3__44,linha8_3__43,linha8_3__42,
              linha8_3__41,linha8_3__40,linha8_3__39,linha8_3__38,linha8_3__37,
              linha8_3__36,linha8_3__35,linha8_3__34,linha8_3__33,linha8_3__32,
              linha8_3__31,linha8_3__30,linha8_3__29,linha8_3__28,linha8_3__27,
              linha8_3__26,linha8_3__25,linha8_3__24,linha8_3__23,linha8_3__22,
              linha8_3__21,linha8_3__20,linha8_3__19,linha8_3__18,linha8_3__17,
              linha8_3__16,linha8_3__15,linha8_3__14,linha8_3__13,linha8_3__12,
              linha8_3__11,linha8_3__10,linha8_3__9,linha8_3__8,linha8_3__7,
              linha8_3__6,linha8_3__5,linha8_3__4,linha8_3__3,linha8_3__2,
              linha8_3__1,linha8_3__0}), .a0 ({linha7_6__63,linha7_6__62,
              linha7_6__61,linha7_6__60,linha7_6__59,linha7_6__58,linha7_6__57,
              linha7_6__56,linha7_6__55,linha7_6__54,linha7_6__53,linha7_6__52,
              linha7_6__51,linha7_6__50,linha7_6__49,linha7_6__48,linha7_6__47,
              linha7_6__46,linha7_6__45,linha7_6__44,linha7_6__43,linha7_6__42,
              linha7_6__41,linha7_6__40,linha7_6__39,linha7_6__38,linha7_6__37,
              linha7_6__36,linha7_6__35,linha7_6__34,linha7_6__33,linha7_6__32,
              linha7_6__31,linha7_6__30,linha7_6__29,linha7_6__28,linha7_6__27,
              linha7_6__26,linha7_6__25,linha7_6__24,linha7_6__23,linha7_6__22,
              linha7_6__21,linha7_6__20,linha7_6__19,linha7_6__18,linha7_6__17,
              linha7_6__16,linha7_6__15,linha7_6__14,linha7_6__13,linha7_6__12,
              linha7_6__11,linha7_6__10,linha7_6__9,linha7_6__8,linha7_6__7,
              linha7_6__6,linha7_6__5,linha7_6__4,linha7_6__3,linha7_6__2,
              linha7_6__1,linha7_6__0}), .s (row_6_rowp_bni4_l)) ;
    Mux2x1_64 row_6_rowp_bni4_muxMin (.r ({y8[63],y8[62],y8[61],y8[60],y8[59],
              y8[58],y8[57],y8[56],y8[55],y8[54],y8[53],y8[52],y8[51],y8[50],
              y8[49],y8[48],y8[47],y8[46],y8[45],y8[44],y8[43],y8[42],y8[41],
              y8[40],y8[39],y8[38],y8[37],y8[36],y8[35],y8[34],y8[33],y8[32],
              y8[31],y8[30],y8[29],y8[28],y8[27],y8[26],y8[25],y8[24],y8[23],
              y8[22],y8[21],y8[20],y8[19],y8[18],y8[17],y8[16],y8[15],y8[14],
              y8[13],y8[12],y8[11],y8[10],y8[9],y8[8],y8[7],y8[6],y8[5],y8[4],
              y8[3],y8[2],y8[1],y8[0]}), .a1 ({linha7_6__63,linha7_6__62,
              linha7_6__61,linha7_6__60,linha7_6__59,linha7_6__58,linha7_6__57,
              linha7_6__56,linha7_6__55,linha7_6__54,linha7_6__53,linha7_6__52,
              linha7_6__51,linha7_6__50,linha7_6__49,linha7_6__48,linha7_6__47,
              linha7_6__46,linha7_6__45,linha7_6__44,linha7_6__43,linha7_6__42,
              linha7_6__41,linha7_6__40,linha7_6__39,linha7_6__38,linha7_6__37,
              linha7_6__36,linha7_6__35,linha7_6__34,linha7_6__33,linha7_6__32,
              linha7_6__31,linha7_6__30,linha7_6__29,linha7_6__28,linha7_6__27,
              linha7_6__26,linha7_6__25,linha7_6__24,linha7_6__23,linha7_6__22,
              linha7_6__21,linha7_6__20,linha7_6__19,linha7_6__18,linha7_6__17,
              linha7_6__16,linha7_6__15,linha7_6__14,linha7_6__13,linha7_6__12,
              linha7_6__11,linha7_6__10,linha7_6__9,linha7_6__8,linha7_6__7,
              linha7_6__6,linha7_6__5,linha7_6__4,linha7_6__3,linha7_6__2,
              linha7_6__1,linha7_6__0}), .a0 ({linha8_3__63,linha8_3__62,
              linha8_3__61,linha8_3__60,linha8_3__59,linha8_3__58,linha8_3__57,
              linha8_3__56,linha8_3__55,linha8_3__54,linha8_3__53,linha8_3__52,
              linha8_3__51,linha8_3__50,linha8_3__49,linha8_3__48,linha8_3__47,
              linha8_3__46,linha8_3__45,linha8_3__44,linha8_3__43,linha8_3__42,
              linha8_3__41,linha8_3__40,linha8_3__39,linha8_3__38,linha8_3__37,
              linha8_3__36,linha8_3__35,linha8_3__34,linha8_3__33,linha8_3__32,
              linha8_3__31,linha8_3__30,linha8_3__29,linha8_3__28,linha8_3__27,
              linha8_3__26,linha8_3__25,linha8_3__24,linha8_3__23,linha8_3__22,
              linha8_3__21,linha8_3__20,linha8_3__19,linha8_3__18,linha8_3__17,
              linha8_3__16,linha8_3__15,linha8_3__14,linha8_3__13,linha8_3__12,
              linha8_3__11,linha8_3__10,linha8_3__9,linha8_3__8,linha8_3__7,
              linha8_3__6,linha8_3__5,linha8_3__4,linha8_3__3,linha8_3__2,
              linha8_3__1,linha8_3__0}), .s (row_6_rowp_bni4_l)) ;
    juntarComparadores_64 row_7_rowi_bni1_Comp (.g (\$dummy [25]), .l (
                          row_7_rowi_bni1_l), .a ({linha2_7__63,linha2_7__62,
                          linha2_7__61,linha2_7__60,linha2_7__59,linha2_7__58,
                          linha2_7__57,linha2_7__56,linha2_7__55,linha2_7__54,
                          linha2_7__53,linha2_7__52,linha2_7__51,linha2_7__50,
                          linha2_7__49,linha2_7__48,linha2_7__47,linha2_7__46,
                          linha2_7__45,linha2_7__44,linha2_7__43,linha2_7__42,
                          linha2_7__41,linha2_7__40,linha2_7__39,linha2_7__38,
                          linha2_7__37,linha2_7__36,linha2_7__35,linha2_7__34,
                          linha2_7__33,linha2_7__32,linha2_7__31,linha2_7__30,
                          linha2_7__29,linha2_7__28,linha2_7__27,linha2_7__26,
                          linha2_7__25,linha2_7__24,linha2_7__23,linha2_7__22,
                          linha2_7__21,linha2_7__20,linha2_7__19,linha2_7__18,
                          linha2_7__17,linha2_7__16,linha2_7__15,linha2_7__14,
                          linha2_7__13,linha2_7__12,linha2_7__11,linha2_7__10,
                          linha2_7__9,linha2_7__8,linha2_7__7,linha2_7__6,
                          linha2_7__5,linha2_7__4,linha2_7__3,linha2_7__2,
                          linha2_7__1,linha2_7__0}), .b ({linha3_7__63,
                          linha3_7__62,linha3_7__61,linha3_7__60,linha3_7__59,
                          linha3_7__58,linha3_7__57,linha3_7__56,linha3_7__55,
                          linha3_7__54,linha3_7__53,linha3_7__52,linha3_7__51,
                          linha3_7__50,linha3_7__49,linha3_7__48,linha3_7__47,
                          linha3_7__46,linha3_7__45,linha3_7__44,linha3_7__43,
                          linha3_7__42,linha3_7__41,linha3_7__40,linha3_7__39,
                          linha3_7__38,linha3_7__37,linha3_7__36,linha3_7__35,
                          linha3_7__34,linha3_7__33,linha3_7__32,linha3_7__31,
                          linha3_7__30,linha3_7__29,linha3_7__28,linha3_7__27,
                          linha3_7__26,linha3_7__25,linha3_7__24,linha3_7__23,
                          linha3_7__22,linha3_7__21,linha3_7__20,linha3_7__19,
                          linha3_7__18,linha3_7__17,linha3_7__16,linha3_7__15,
                          linha3_7__14,linha3_7__13,linha3_7__12,linha3_7__11,
                          linha3_7__10,linha3_7__9,linha3_7__8,linha3_7__7,
                          linha3_7__6,linha3_7__5,linha3_7__4,linha3_7__3,
                          linha3_7__2,linha3_7__1,linha3_7__0})) ;
    Mux2x1_64 row_7_rowi_bni1_muxMax (.r ({y2[63],y2[62],y2[61],y2[60],y2[59],
              y2[58],y2[57],y2[56],y2[55],y2[54],y2[53],y2[52],y2[51],y2[50],
              y2[49],y2[48],y2[47],y2[46],y2[45],y2[44],y2[43],y2[42],y2[41],
              y2[40],y2[39],y2[38],y2[37],y2[36],y2[35],y2[34],y2[33],y2[32],
              y2[31],y2[30],y2[29],y2[28],y2[27],y2[26],y2[25],y2[24],y2[23],
              y2[22],y2[21],y2[20],y2[19],y2[18],y2[17],y2[16],y2[15],y2[14],
              y2[13],y2[12],y2[11],y2[10],y2[9],y2[8],y2[7],y2[6],y2[5],y2[4],
              y2[3],y2[2],y2[1],y2[0]}), .a1 ({linha3_7__63,linha3_7__62,
              linha3_7__61,linha3_7__60,linha3_7__59,linha3_7__58,linha3_7__57,
              linha3_7__56,linha3_7__55,linha3_7__54,linha3_7__53,linha3_7__52,
              linha3_7__51,linha3_7__50,linha3_7__49,linha3_7__48,linha3_7__47,
              linha3_7__46,linha3_7__45,linha3_7__44,linha3_7__43,linha3_7__42,
              linha3_7__41,linha3_7__40,linha3_7__39,linha3_7__38,linha3_7__37,
              linha3_7__36,linha3_7__35,linha3_7__34,linha3_7__33,linha3_7__32,
              linha3_7__31,linha3_7__30,linha3_7__29,linha3_7__28,linha3_7__27,
              linha3_7__26,linha3_7__25,linha3_7__24,linha3_7__23,linha3_7__22,
              linha3_7__21,linha3_7__20,linha3_7__19,linha3_7__18,linha3_7__17,
              linha3_7__16,linha3_7__15,linha3_7__14,linha3_7__13,linha3_7__12,
              linha3_7__11,linha3_7__10,linha3_7__9,linha3_7__8,linha3_7__7,
              linha3_7__6,linha3_7__5,linha3_7__4,linha3_7__3,linha3_7__2,
              linha3_7__1,linha3_7__0}), .a0 ({linha2_7__63,linha2_7__62,
              linha2_7__61,linha2_7__60,linha2_7__59,linha2_7__58,linha2_7__57,
              linha2_7__56,linha2_7__55,linha2_7__54,linha2_7__53,linha2_7__52,
              linha2_7__51,linha2_7__50,linha2_7__49,linha2_7__48,linha2_7__47,
              linha2_7__46,linha2_7__45,linha2_7__44,linha2_7__43,linha2_7__42,
              linha2_7__41,linha2_7__40,linha2_7__39,linha2_7__38,linha2_7__37,
              linha2_7__36,linha2_7__35,linha2_7__34,linha2_7__33,linha2_7__32,
              linha2_7__31,linha2_7__30,linha2_7__29,linha2_7__28,linha2_7__27,
              linha2_7__26,linha2_7__25,linha2_7__24,linha2_7__23,linha2_7__22,
              linha2_7__21,linha2_7__20,linha2_7__19,linha2_7__18,linha2_7__17,
              linha2_7__16,linha2_7__15,linha2_7__14,linha2_7__13,linha2_7__12,
              linha2_7__11,linha2_7__10,linha2_7__9,linha2_7__8,linha2_7__7,
              linha2_7__6,linha2_7__5,linha2_7__4,linha2_7__3,linha2_7__2,
              linha2_7__1,linha2_7__0}), .s (row_7_rowi_bni1_l)) ;
    Mux2x1_64 row_7_rowi_bni1_muxMin (.r ({y3[63],y3[62],y3[61],y3[60],y3[59],
              y3[58],y3[57],y3[56],y3[55],y3[54],y3[53],y3[52],y3[51],y3[50],
              y3[49],y3[48],y3[47],y3[46],y3[45],y3[44],y3[43],y3[42],y3[41],
              y3[40],y3[39],y3[38],y3[37],y3[36],y3[35],y3[34],y3[33],y3[32],
              y3[31],y3[30],y3[29],y3[28],y3[27],y3[26],y3[25],y3[24],y3[23],
              y3[22],y3[21],y3[20],y3[19],y3[18],y3[17],y3[16],y3[15],y3[14],
              y3[13],y3[12],y3[11],y3[10],y3[9],y3[8],y3[7],y3[6],y3[5],y3[4],
              y3[3],y3[2],y3[1],y3[0]}), .a1 ({linha2_7__63,linha2_7__62,
              linha2_7__61,linha2_7__60,linha2_7__59,linha2_7__58,linha2_7__57,
              linha2_7__56,linha2_7__55,linha2_7__54,linha2_7__53,linha2_7__52,
              linha2_7__51,linha2_7__50,linha2_7__49,linha2_7__48,linha2_7__47,
              linha2_7__46,linha2_7__45,linha2_7__44,linha2_7__43,linha2_7__42,
              linha2_7__41,linha2_7__40,linha2_7__39,linha2_7__38,linha2_7__37,
              linha2_7__36,linha2_7__35,linha2_7__34,linha2_7__33,linha2_7__32,
              linha2_7__31,linha2_7__30,linha2_7__29,linha2_7__28,linha2_7__27,
              linha2_7__26,linha2_7__25,linha2_7__24,linha2_7__23,linha2_7__22,
              linha2_7__21,linha2_7__20,linha2_7__19,linha2_7__18,linha2_7__17,
              linha2_7__16,linha2_7__15,linha2_7__14,linha2_7__13,linha2_7__12,
              linha2_7__11,linha2_7__10,linha2_7__9,linha2_7__8,linha2_7__7,
              linha2_7__6,linha2_7__5,linha2_7__4,linha2_7__3,linha2_7__2,
              linha2_7__1,linha2_7__0}), .a0 ({linha3_7__63,linha3_7__62,
              linha3_7__61,linha3_7__60,linha3_7__59,linha3_7__58,linha3_7__57,
              linha3_7__56,linha3_7__55,linha3_7__54,linha3_7__53,linha3_7__52,
              linha3_7__51,linha3_7__50,linha3_7__49,linha3_7__48,linha3_7__47,
              linha3_7__46,linha3_7__45,linha3_7__44,linha3_7__43,linha3_7__42,
              linha3_7__41,linha3_7__40,linha3_7__39,linha3_7__38,linha3_7__37,
              linha3_7__36,linha3_7__35,linha3_7__34,linha3_7__33,linha3_7__32,
              linha3_7__31,linha3_7__30,linha3_7__29,linha3_7__28,linha3_7__27,
              linha3_7__26,linha3_7__25,linha3_7__24,linha3_7__23,linha3_7__22,
              linha3_7__21,linha3_7__20,linha3_7__19,linha3_7__18,linha3_7__17,
              linha3_7__16,linha3_7__15,linha3_7__14,linha3_7__13,linha3_7__12,
              linha3_7__11,linha3_7__10,linha3_7__9,linha3_7__8,linha3_7__7,
              linha3_7__6,linha3_7__5,linha3_7__4,linha3_7__3,linha3_7__2,
              linha3_7__1,linha3_7__0}), .s (row_7_rowi_bni1_l)) ;
    juntarComparadores_64 row_7_rowi_bni2_Comp (.g (\$dummy [26]), .l (
                          row_7_rowi_bni2_l), .a ({linha4_7__63,linha4_7__62,
                          linha4_7__61,linha4_7__60,linha4_7__59,linha4_7__58,
                          linha4_7__57,linha4_7__56,linha4_7__55,linha4_7__54,
                          linha4_7__53,linha4_7__52,linha4_7__51,linha4_7__50,
                          linha4_7__49,linha4_7__48,linha4_7__47,linha4_7__46,
                          linha4_7__45,linha4_7__44,linha4_7__43,linha4_7__42,
                          linha4_7__41,linha4_7__40,linha4_7__39,linha4_7__38,
                          linha4_7__37,linha4_7__36,linha4_7__35,linha4_7__34,
                          linha4_7__33,linha4_7__32,linha4_7__31,linha4_7__30,
                          linha4_7__29,linha4_7__28,linha4_7__27,linha4_7__26,
                          linha4_7__25,linha4_7__24,linha4_7__23,linha4_7__22,
                          linha4_7__21,linha4_7__20,linha4_7__19,linha4_7__18,
                          linha4_7__17,linha4_7__16,linha4_7__15,linha4_7__14,
                          linha4_7__13,linha4_7__12,linha4_7__11,linha4_7__10,
                          linha4_7__9,linha4_7__8,linha4_7__7,linha4_7__6,
                          linha4_7__5,linha4_7__4,linha4_7__3,linha4_7__2,
                          linha4_7__1,linha4_7__0}), .b ({linha5_7__63,
                          linha5_7__62,linha5_7__61,linha5_7__60,linha5_7__59,
                          linha5_7__58,linha5_7__57,linha5_7__56,linha5_7__55,
                          linha5_7__54,linha5_7__53,linha5_7__52,linha5_7__51,
                          linha5_7__50,linha5_7__49,linha5_7__48,linha5_7__47,
                          linha5_7__46,linha5_7__45,linha5_7__44,linha5_7__43,
                          linha5_7__42,linha5_7__41,linha5_7__40,linha5_7__39,
                          linha5_7__38,linha5_7__37,linha5_7__36,linha5_7__35,
                          linha5_7__34,linha5_7__33,linha5_7__32,linha5_7__31,
                          linha5_7__30,linha5_7__29,linha5_7__28,linha5_7__27,
                          linha5_7__26,linha5_7__25,linha5_7__24,linha5_7__23,
                          linha5_7__22,linha5_7__21,linha5_7__20,linha5_7__19,
                          linha5_7__18,linha5_7__17,linha5_7__16,linha5_7__15,
                          linha5_7__14,linha5_7__13,linha5_7__12,linha5_7__11,
                          linha5_7__10,linha5_7__9,linha5_7__8,linha5_7__7,
                          linha5_7__6,linha5_7__5,linha5_7__4,linha5_7__3,
                          linha5_7__2,linha5_7__1,linha5_7__0})) ;
    Mux2x1_64 row_7_rowi_bni2_muxMax (.r ({y4[63],y4[62],y4[61],y4[60],y4[59],
              y4[58],y4[57],y4[56],y4[55],y4[54],y4[53],y4[52],y4[51],y4[50],
              y4[49],y4[48],y4[47],y4[46],y4[45],y4[44],y4[43],y4[42],y4[41],
              y4[40],y4[39],y4[38],y4[37],y4[36],y4[35],y4[34],y4[33],y4[32],
              y4[31],y4[30],y4[29],y4[28],y4[27],y4[26],y4[25],y4[24],y4[23],
              y4[22],y4[21],y4[20],y4[19],y4[18],y4[17],y4[16],y4[15],y4[14],
              y4[13],y4[12],y4[11],y4[10],y4[9],y4[8],y4[7],y4[6],y4[5],y4[4],
              y4[3],y4[2],y4[1],y4[0]}), .a1 ({linha5_7__63,linha5_7__62,
              linha5_7__61,linha5_7__60,linha5_7__59,linha5_7__58,linha5_7__57,
              linha5_7__56,linha5_7__55,linha5_7__54,linha5_7__53,linha5_7__52,
              linha5_7__51,linha5_7__50,linha5_7__49,linha5_7__48,linha5_7__47,
              linha5_7__46,linha5_7__45,linha5_7__44,linha5_7__43,linha5_7__42,
              linha5_7__41,linha5_7__40,linha5_7__39,linha5_7__38,linha5_7__37,
              linha5_7__36,linha5_7__35,linha5_7__34,linha5_7__33,linha5_7__32,
              linha5_7__31,linha5_7__30,linha5_7__29,linha5_7__28,linha5_7__27,
              linha5_7__26,linha5_7__25,linha5_7__24,linha5_7__23,linha5_7__22,
              linha5_7__21,linha5_7__20,linha5_7__19,linha5_7__18,linha5_7__17,
              linha5_7__16,linha5_7__15,linha5_7__14,linha5_7__13,linha5_7__12,
              linha5_7__11,linha5_7__10,linha5_7__9,linha5_7__8,linha5_7__7,
              linha5_7__6,linha5_7__5,linha5_7__4,linha5_7__3,linha5_7__2,
              linha5_7__1,linha5_7__0}), .a0 ({linha4_7__63,linha4_7__62,
              linha4_7__61,linha4_7__60,linha4_7__59,linha4_7__58,linha4_7__57,
              linha4_7__56,linha4_7__55,linha4_7__54,linha4_7__53,linha4_7__52,
              linha4_7__51,linha4_7__50,linha4_7__49,linha4_7__48,linha4_7__47,
              linha4_7__46,linha4_7__45,linha4_7__44,linha4_7__43,linha4_7__42,
              linha4_7__41,linha4_7__40,linha4_7__39,linha4_7__38,linha4_7__37,
              linha4_7__36,linha4_7__35,linha4_7__34,linha4_7__33,linha4_7__32,
              linha4_7__31,linha4_7__30,linha4_7__29,linha4_7__28,linha4_7__27,
              linha4_7__26,linha4_7__25,linha4_7__24,linha4_7__23,linha4_7__22,
              linha4_7__21,linha4_7__20,linha4_7__19,linha4_7__18,linha4_7__17,
              linha4_7__16,linha4_7__15,linha4_7__14,linha4_7__13,linha4_7__12,
              linha4_7__11,linha4_7__10,linha4_7__9,linha4_7__8,linha4_7__7,
              linha4_7__6,linha4_7__5,linha4_7__4,linha4_7__3,linha4_7__2,
              linha4_7__1,linha4_7__0}), .s (row_7_rowi_bni2_l)) ;
    Mux2x1_64 row_7_rowi_bni2_muxMin (.r ({y5[63],y5[62],y5[61],y5[60],y5[59],
              y5[58],y5[57],y5[56],y5[55],y5[54],y5[53],y5[52],y5[51],y5[50],
              y5[49],y5[48],y5[47],y5[46],y5[45],y5[44],y5[43],y5[42],y5[41],
              y5[40],y5[39],y5[38],y5[37],y5[36],y5[35],y5[34],y5[33],y5[32],
              y5[31],y5[30],y5[29],y5[28],y5[27],y5[26],y5[25],y5[24],y5[23],
              y5[22],y5[21],y5[20],y5[19],y5[18],y5[17],y5[16],y5[15],y5[14],
              y5[13],y5[12],y5[11],y5[10],y5[9],y5[8],y5[7],y5[6],y5[5],y5[4],
              y5[3],y5[2],y5[1],y5[0]}), .a1 ({linha4_7__63,linha4_7__62,
              linha4_7__61,linha4_7__60,linha4_7__59,linha4_7__58,linha4_7__57,
              linha4_7__56,linha4_7__55,linha4_7__54,linha4_7__53,linha4_7__52,
              linha4_7__51,linha4_7__50,linha4_7__49,linha4_7__48,linha4_7__47,
              linha4_7__46,linha4_7__45,linha4_7__44,linha4_7__43,linha4_7__42,
              linha4_7__41,linha4_7__40,linha4_7__39,linha4_7__38,linha4_7__37,
              linha4_7__36,linha4_7__35,linha4_7__34,linha4_7__33,linha4_7__32,
              linha4_7__31,linha4_7__30,linha4_7__29,linha4_7__28,linha4_7__27,
              linha4_7__26,linha4_7__25,linha4_7__24,linha4_7__23,linha4_7__22,
              linha4_7__21,linha4_7__20,linha4_7__19,linha4_7__18,linha4_7__17,
              linha4_7__16,linha4_7__15,linha4_7__14,linha4_7__13,linha4_7__12,
              linha4_7__11,linha4_7__10,linha4_7__9,linha4_7__8,linha4_7__7,
              linha4_7__6,linha4_7__5,linha4_7__4,linha4_7__3,linha4_7__2,
              linha4_7__1,linha4_7__0}), .a0 ({linha5_7__63,linha5_7__62,
              linha5_7__61,linha5_7__60,linha5_7__59,linha5_7__58,linha5_7__57,
              linha5_7__56,linha5_7__55,linha5_7__54,linha5_7__53,linha5_7__52,
              linha5_7__51,linha5_7__50,linha5_7__49,linha5_7__48,linha5_7__47,
              linha5_7__46,linha5_7__45,linha5_7__44,linha5_7__43,linha5_7__42,
              linha5_7__41,linha5_7__40,linha5_7__39,linha5_7__38,linha5_7__37,
              linha5_7__36,linha5_7__35,linha5_7__34,linha5_7__33,linha5_7__32,
              linha5_7__31,linha5_7__30,linha5_7__29,linha5_7__28,linha5_7__27,
              linha5_7__26,linha5_7__25,linha5_7__24,linha5_7__23,linha5_7__22,
              linha5_7__21,linha5_7__20,linha5_7__19,linha5_7__18,linha5_7__17,
              linha5_7__16,linha5_7__15,linha5_7__14,linha5_7__13,linha5_7__12,
              linha5_7__11,linha5_7__10,linha5_7__9,linha5_7__8,linha5_7__7,
              linha5_7__6,linha5_7__5,linha5_7__4,linha5_7__3,linha5_7__2,
              linha5_7__1,linha5_7__0}), .s (row_7_rowi_bni2_l)) ;
    juntarComparadores_64 row_7_rowi_bni3_Comp (.g (\$dummy [27]), .l (
                          row_7_rowi_bni3_l), .a ({linha6_7__63,linha6_7__62,
                          linha6_7__61,linha6_7__60,linha6_7__59,linha6_7__58,
                          linha6_7__57,linha6_7__56,linha6_7__55,linha6_7__54,
                          linha6_7__53,linha6_7__52,linha6_7__51,linha6_7__50,
                          linha6_7__49,linha6_7__48,linha6_7__47,linha6_7__46,
                          linha6_7__45,linha6_7__44,linha6_7__43,linha6_7__42,
                          linha6_7__41,linha6_7__40,linha6_7__39,linha6_7__38,
                          linha6_7__37,linha6_7__36,linha6_7__35,linha6_7__34,
                          linha6_7__33,linha6_7__32,linha6_7__31,linha6_7__30,
                          linha6_7__29,linha6_7__28,linha6_7__27,linha6_7__26,
                          linha6_7__25,linha6_7__24,linha6_7__23,linha6_7__22,
                          linha6_7__21,linha6_7__20,linha6_7__19,linha6_7__18,
                          linha6_7__17,linha6_7__16,linha6_7__15,linha6_7__14,
                          linha6_7__13,linha6_7__12,linha6_7__11,linha6_7__10,
                          linha6_7__9,linha6_7__8,linha6_7__7,linha6_7__6,
                          linha6_7__5,linha6_7__4,linha6_7__3,linha6_7__2,
                          linha6_7__1,linha6_7__0}), .b ({linha7_7__63,
                          linha7_7__62,linha7_7__61,linha7_7__60,linha7_7__59,
                          linha7_7__58,linha7_7__57,linha7_7__56,linha7_7__55,
                          linha7_7__54,linha7_7__53,linha7_7__52,linha7_7__51,
                          linha7_7__50,linha7_7__49,linha7_7__48,linha7_7__47,
                          linha7_7__46,linha7_7__45,linha7_7__44,linha7_7__43,
                          linha7_7__42,linha7_7__41,linha7_7__40,linha7_7__39,
                          linha7_7__38,linha7_7__37,linha7_7__36,linha7_7__35,
                          linha7_7__34,linha7_7__33,linha7_7__32,linha7_7__31,
                          linha7_7__30,linha7_7__29,linha7_7__28,linha7_7__27,
                          linha7_7__26,linha7_7__25,linha7_7__24,linha7_7__23,
                          linha7_7__22,linha7_7__21,linha7_7__20,linha7_7__19,
                          linha7_7__18,linha7_7__17,linha7_7__16,linha7_7__15,
                          linha7_7__14,linha7_7__13,linha7_7__12,linha7_7__11,
                          linha7_7__10,linha7_7__9,linha7_7__8,linha7_7__7,
                          linha7_7__6,linha7_7__5,linha7_7__4,linha7_7__3,
                          linha7_7__2,linha7_7__1,linha7_7__0})) ;
    Mux2x1_64 row_7_rowi_bni3_muxMax (.r ({y6[63],y6[62],y6[61],y6[60],y6[59],
              y6[58],y6[57],y6[56],y6[55],y6[54],y6[53],y6[52],y6[51],y6[50],
              y6[49],y6[48],y6[47],y6[46],y6[45],y6[44],y6[43],y6[42],y6[41],
              y6[40],y6[39],y6[38],y6[37],y6[36],y6[35],y6[34],y6[33],y6[32],
              y6[31],y6[30],y6[29],y6[28],y6[27],y6[26],y6[25],y6[24],y6[23],
              y6[22],y6[21],y6[20],y6[19],y6[18],y6[17],y6[16],y6[15],y6[14],
              y6[13],y6[12],y6[11],y6[10],y6[9],y6[8],y6[7],y6[6],y6[5],y6[4],
              y6[3],y6[2],y6[1],y6[0]}), .a1 ({linha7_7__63,linha7_7__62,
              linha7_7__61,linha7_7__60,linha7_7__59,linha7_7__58,linha7_7__57,
              linha7_7__56,linha7_7__55,linha7_7__54,linha7_7__53,linha7_7__52,
              linha7_7__51,linha7_7__50,linha7_7__49,linha7_7__48,linha7_7__47,
              linha7_7__46,linha7_7__45,linha7_7__44,linha7_7__43,linha7_7__42,
              linha7_7__41,linha7_7__40,linha7_7__39,linha7_7__38,linha7_7__37,
              linha7_7__36,linha7_7__35,linha7_7__34,linha7_7__33,linha7_7__32,
              linha7_7__31,linha7_7__30,linha7_7__29,linha7_7__28,linha7_7__27,
              linha7_7__26,linha7_7__25,linha7_7__24,linha7_7__23,linha7_7__22,
              linha7_7__21,linha7_7__20,linha7_7__19,linha7_7__18,linha7_7__17,
              linha7_7__16,linha7_7__15,linha7_7__14,linha7_7__13,linha7_7__12,
              linha7_7__11,linha7_7__10,linha7_7__9,linha7_7__8,linha7_7__7,
              linha7_7__6,linha7_7__5,linha7_7__4,linha7_7__3,linha7_7__2,
              linha7_7__1,linha7_7__0}), .a0 ({linha6_7__63,linha6_7__62,
              linha6_7__61,linha6_7__60,linha6_7__59,linha6_7__58,linha6_7__57,
              linha6_7__56,linha6_7__55,linha6_7__54,linha6_7__53,linha6_7__52,
              linha6_7__51,linha6_7__50,linha6_7__49,linha6_7__48,linha6_7__47,
              linha6_7__46,linha6_7__45,linha6_7__44,linha6_7__43,linha6_7__42,
              linha6_7__41,linha6_7__40,linha6_7__39,linha6_7__38,linha6_7__37,
              linha6_7__36,linha6_7__35,linha6_7__34,linha6_7__33,linha6_7__32,
              linha6_7__31,linha6_7__30,linha6_7__29,linha6_7__28,linha6_7__27,
              linha6_7__26,linha6_7__25,linha6_7__24,linha6_7__23,linha6_7__22,
              linha6_7__21,linha6_7__20,linha6_7__19,linha6_7__18,linha6_7__17,
              linha6_7__16,linha6_7__15,linha6_7__14,linha6_7__13,linha6_7__12,
              linha6_7__11,linha6_7__10,linha6_7__9,linha6_7__8,linha6_7__7,
              linha6_7__6,linha6_7__5,linha6_7__4,linha6_7__3,linha6_7__2,
              linha6_7__1,linha6_7__0}), .s (row_7_rowi_bni3_l)) ;
    Mux2x1_64 row_7_rowi_bni3_muxMin (.r ({y7[63],y7[62],y7[61],y7[60],y7[59],
              y7[58],y7[57],y7[56],y7[55],y7[54],y7[53],y7[52],y7[51],y7[50],
              y7[49],y7[48],y7[47],y7[46],y7[45],y7[44],y7[43],y7[42],y7[41],
              y7[40],y7[39],y7[38],y7[37],y7[36],y7[35],y7[34],y7[33],y7[32],
              y7[31],y7[30],y7[29],y7[28],y7[27],y7[26],y7[25],y7[24],y7[23],
              y7[22],y7[21],y7[20],y7[19],y7[18],y7[17],y7[16],y7[15],y7[14],
              y7[13],y7[12],y7[11],y7[10],y7[9],y7[8],y7[7],y7[6],y7[5],y7[4],
              y7[3],y7[2],y7[1],y7[0]}), .a1 ({linha6_7__63,linha6_7__62,
              linha6_7__61,linha6_7__60,linha6_7__59,linha6_7__58,linha6_7__57,
              linha6_7__56,linha6_7__55,linha6_7__54,linha6_7__53,linha6_7__52,
              linha6_7__51,linha6_7__50,linha6_7__49,linha6_7__48,linha6_7__47,
              linha6_7__46,linha6_7__45,linha6_7__44,linha6_7__43,linha6_7__42,
              linha6_7__41,linha6_7__40,linha6_7__39,linha6_7__38,linha6_7__37,
              linha6_7__36,linha6_7__35,linha6_7__34,linha6_7__33,linha6_7__32,
              linha6_7__31,linha6_7__30,linha6_7__29,linha6_7__28,linha6_7__27,
              linha6_7__26,linha6_7__25,linha6_7__24,linha6_7__23,linha6_7__22,
              linha6_7__21,linha6_7__20,linha6_7__19,linha6_7__18,linha6_7__17,
              linha6_7__16,linha6_7__15,linha6_7__14,linha6_7__13,linha6_7__12,
              linha6_7__11,linha6_7__10,linha6_7__9,linha6_7__8,linha6_7__7,
              linha6_7__6,linha6_7__5,linha6_7__4,linha6_7__3,linha6_7__2,
              linha6_7__1,linha6_7__0}), .a0 ({linha7_7__63,linha7_7__62,
              linha7_7__61,linha7_7__60,linha7_7__59,linha7_7__58,linha7_7__57,
              linha7_7__56,linha7_7__55,linha7_7__54,linha7_7__53,linha7_7__52,
              linha7_7__51,linha7_7__50,linha7_7__49,linha7_7__48,linha7_7__47,
              linha7_7__46,linha7_7__45,linha7_7__44,linha7_7__43,linha7_7__42,
              linha7_7__41,linha7_7__40,linha7_7__39,linha7_7__38,linha7_7__37,
              linha7_7__36,linha7_7__35,linha7_7__34,linha7_7__33,linha7_7__32,
              linha7_7__31,linha7_7__30,linha7_7__29,linha7_7__28,linha7_7__27,
              linha7_7__26,linha7_7__25,linha7_7__24,linha7_7__23,linha7_7__22,
              linha7_7__21,linha7_7__20,linha7_7__19,linha7_7__18,linha7_7__17,
              linha7_7__16,linha7_7__15,linha7_7__14,linha7_7__13,linha7_7__12,
              linha7_7__11,linha7_7__10,linha7_7__9,linha7_7__8,linha7_7__7,
              linha7_7__6,linha7_7__5,linha7_7__4,linha7_7__3,linha7_7__2,
              linha7_7__1,linha7_7__0}), .s (row_7_rowi_bni3_l)) ;
    AN1T0 ix8126 (.X (nx8127), .A (row_0_rowp_bni1_l)) ;
endmodule


module AN1T0 ( X, A ) ;

    output X ;
    input A ;




    assign X = A ;
endmodule


module Mux2x1_64 ( r, a1, a0, s ) ;

    output [63:0]r ;
    input [63:0]a1 ;
    input [63:0]a0 ;
    input s ;

    wire nx639, nx641;



    MX2T0 ix7 (.X (r[0]), .A (a1[0]), .B (a0[0]), .S (nx639)) ;
    MX2T0 ix15 (.X (r[1]), .A (a1[1]), .B (a0[1]), .S (nx639)) ;
    MX2T0 ix23 (.X (r[2]), .A (a1[2]), .B (a0[2]), .S (nx639)) ;
    MX2T0 ix31 (.X (r[3]), .A (a1[3]), .B (a0[3]), .S (nx639)) ;
    MX2T0 ix39 (.X (r[4]), .A (a1[4]), .B (a0[4]), .S (nx639)) ;
    MX2T0 ix47 (.X (r[5]), .A (a1[5]), .B (a0[5]), .S (nx639)) ;
    MX2T0 ix55 (.X (r[6]), .A (a1[6]), .B (a0[6]), .S (nx639)) ;
    MX2T0 ix63 (.X (r[7]), .A (a1[7]), .B (a0[7]), .S (nx639)) ;
    MX2T0 ix71 (.X (r[8]), .A (a1[8]), .B (a0[8]), .S (nx639)) ;
    MX2T0 ix79 (.X (r[9]), .A (a1[9]), .B (a0[9]), .S (nx639)) ;
    MX2T0 ix87 (.X (r[10]), .A (a1[10]), .B (a0[10]), .S (nx639)) ;
    MX2T0 ix95 (.X (r[11]), .A (a1[11]), .B (a0[11]), .S (nx639)) ;
    MX2T0 ix103 (.X (r[12]), .A (a1[12]), .B (a0[12]), .S (nx639)) ;
    MX2T0 ix111 (.X (r[13]), .A (a1[13]), .B (a0[13]), .S (nx639)) ;
    MX2T0 ix119 (.X (r[14]), .A (a1[14]), .B (a0[14]), .S (nx639)) ;
    MX2T0 ix127 (.X (r[15]), .A (a1[15]), .B (a0[15]), .S (nx639)) ;
    MX2T0 ix135 (.X (r[16]), .A (a1[16]), .B (a0[16]), .S (nx639)) ;
    MX2T0 ix143 (.X (r[17]), .A (a1[17]), .B (a0[17]), .S (nx639)) ;
    MX2T0 ix151 (.X (r[18]), .A (a1[18]), .B (a0[18]), .S (nx639)) ;
    MX2T0 ix159 (.X (r[19]), .A (a1[19]), .B (a0[19]), .S (nx639)) ;
    MX2T0 ix167 (.X (r[20]), .A (a1[20]), .B (a0[20]), .S (nx639)) ;
    MX2T0 ix175 (.X (r[21]), .A (a1[21]), .B (a0[21]), .S (nx639)) ;
    MX2T0 ix183 (.X (r[22]), .A (a1[22]), .B (a0[22]), .S (nx639)) ;
    MX2T0 ix191 (.X (r[23]), .A (a1[23]), .B (a0[23]), .S (nx639)) ;
    MX2T0 ix199 (.X (r[24]), .A (a1[24]), .B (a0[24]), .S (nx639)) ;
    MX2T0 ix207 (.X (r[25]), .A (a1[25]), .B (a0[25]), .S (nx639)) ;
    MX2T0 ix215 (.X (r[26]), .A (a1[26]), .B (a0[26]), .S (nx639)) ;
    MX2T0 ix223 (.X (r[27]), .A (a1[27]), .B (a0[27]), .S (nx639)) ;
    MX2T0 ix231 (.X (r[28]), .A (a1[28]), .B (a0[28]), .S (nx639)) ;
    MX2T0 ix239 (.X (r[29]), .A (a1[29]), .B (a0[29]), .S (nx639)) ;
    MX2T0 ix247 (.X (r[30]), .A (a1[30]), .B (a0[30]), .S (nx639)) ;
    MX2T0 ix255 (.X (r[31]), .A (a1[31]), .B (a0[31]), .S (nx639)) ;
    MX2T0 ix263 (.X (r[32]), .A (a1[32]), .B (a0[32]), .S (nx639)) ;
    MX2T0 ix271 (.X (r[33]), .A (a1[33]), .B (a0[33]), .S (nx639)) ;
    MX2T0 ix279 (.X (r[34]), .A (a1[34]), .B (a0[34]), .S (nx639)) ;
    MX2T0 ix287 (.X (r[35]), .A (a1[35]), .B (a0[35]), .S (nx639)) ;
    MX2T0 ix295 (.X (r[36]), .A (a1[36]), .B (a0[36]), .S (nx639)) ;
    MX2T0 ix303 (.X (r[37]), .A (a1[37]), .B (a0[37]), .S (nx639)) ;
    MX2T0 ix311 (.X (r[38]), .A (a1[38]), .B (a0[38]), .S (nx639)) ;
    MX2T0 ix319 (.X (r[39]), .A (a1[39]), .B (a0[39]), .S (nx639)) ;
    MX2T0 ix327 (.X (r[40]), .A (a1[40]), .B (a0[40]), .S (nx639)) ;
    MX2T0 ix335 (.X (r[41]), .A (a1[41]), .B (a0[41]), .S (nx639)) ;
    MX2T0 ix343 (.X (r[42]), .A (a1[42]), .B (a0[42]), .S (nx641)) ;
    MX2T0 ix351 (.X (r[43]), .A (a1[43]), .B (a0[43]), .S (nx641)) ;
    MX2T0 ix359 (.X (r[44]), .A (a1[44]), .B (a0[44]), .S (nx641)) ;
    MX2T0 ix367 (.X (r[45]), .A (a1[45]), .B (a0[45]), .S (nx641)) ;
    MX2T0 ix375 (.X (r[46]), .A (a1[46]), .B (a0[46]), .S (nx641)) ;
    MX2T0 ix383 (.X (r[47]), .A (a1[47]), .B (a0[47]), .S (nx641)) ;
    MX2T0 ix391 (.X (r[48]), .A (a1[48]), .B (a0[48]), .S (nx641)) ;
    MX2T0 ix399 (.X (r[49]), .A (a1[49]), .B (a0[49]), .S (nx641)) ;
    MX2T0 ix407 (.X (r[50]), .A (a1[50]), .B (a0[50]), .S (nx641)) ;
    MX2T0 ix415 (.X (r[51]), .A (a1[51]), .B (a0[51]), .S (nx641)) ;
    MX2T0 ix423 (.X (r[52]), .A (a1[52]), .B (a0[52]), .S (nx641)) ;
    MX2T0 ix431 (.X (r[53]), .A (a1[53]), .B (a0[53]), .S (nx641)) ;
    MX2T0 ix439 (.X (r[54]), .A (a1[54]), .B (a0[54]), .S (nx641)) ;
    MX2T0 ix447 (.X (r[55]), .A (a1[55]), .B (a0[55]), .S (nx641)) ;
    MX2T0 ix455 (.X (r[56]), .A (a1[56]), .B (a0[56]), .S (nx641)) ;
    MX2T0 ix463 (.X (r[57]), .A (a1[57]), .B (a0[57]), .S (nx641)) ;
    MX2T0 ix471 (.X (r[58]), .A (a1[58]), .B (a0[58]), .S (nx641)) ;
    MX2T0 ix479 (.X (r[59]), .A (a1[59]), .B (a0[59]), .S (nx641)) ;
    MX2T0 ix487 (.X (r[60]), .A (a1[60]), .B (a0[60]), .S (nx641)) ;
    MX2T0 ix495 (.X (r[61]), .A (a1[61]), .B (a0[61]), .S (nx641)) ;
    MX2T0 ix503 (.X (r[62]), .A (a1[62]), .B (a0[62]), .S (nx641)) ;
    MX2T0 ix511 (.X (r[63]), .A (a1[63]), .B (a0[63]), .S (nx641)) ;
    AN1V1 ix638 (.X (nx639), .A (s)) ;
    AN1V1 ix640 (.X (nx641), .A (s)) ;
endmodule


module AN1V1 ( X, A ) ;

    output X ;
    input A ;




    assign X = A ;
endmodule


module MX2T0 ( X, A, B, S ) ;

    output X ;
    input A ;
    input B ;
    input S ;

    wire NOT_S, nx2, nx4;



    assign NOT_S = ~S ;
    and (nx2, B, NOT_S) ;
    and (nx4, A, S) ;
    or (X, nx2, nx4) ;
endmodule


module juntarComparadores_64 ( g, l, a, b ) ;

    output g ;
    output l ;
    input [63:0]a ;
    input [63:0]b ;

    wire nx28, nx48, nx58, nx88, nx98, nx128, nx138, nx168, nx178, nx208, nx218, 
         nx248, nx258, nx288, nx298, nx328, nx338, nx368, nx378, nx408, nx418, 
         nx448, nx458, nx488, nx498, nx528, nx538, nx568, nx578, nx608, nx618, 
         nx648, nx658, nx688, nx698, nx728, nx738, nx768, nx778, nx808, nx818, 
         nx848, nx858, nx888, nx898, nx928, nx938, nx968, nx978, nx1008, nx1018, 
         nx1048, nx1058, nx1088, nx1098, nx1128, nx1138, nx1168, nx1178, nx1208, 
         nx1218, nx1238, nx1248, nx939, nx941, nx943, nx945, nx947, nx949, nx951, 
         nx953, nx955, nx957, nx959, nx961, nx963, nx965, nx967, nx969, nx971, 
         nx973, nx975, nx977, nx979, nx981, nx983, nx985, nx987, nx989, nx991, 
         nx993, nx995, nx997, nx999, nx1001, nx1003, nx1005, nx1007, nx1009, 
         nx1011, nx1013, nx1015, nx1017, nx1019, nx1021, nx1023, nx1025, nx1027, 
         nx1029, nx1031, nx1033, nx1035, nx1037, nx1039, nx1041, nx1043, nx1045, 
         nx1047, nx1049, nx1051, nx1053, nx1055, nx1057, nx1059, nx1061, nx1063, 
         nx1065, nx1067, nx1069, nx1071, nx1073, nx1075, nx1077, nx1079, nx1081, 
         nx1083, nx1085, nx1087, nx1089, nx1091, nx1093, nx1095, nx1097, nx1099, 
         nx1101, nx1103, nx1105, nx1107, nx1109, nx1111, nx1113, nx1115, nx1117, 
         nx1119, nx1121, nx1123, nx1125, nx1127, nx1129, nx1131, nx1133, nx1135, 
         nx1137, nx1139, nx1141, nx1143, nx1145, nx1147, nx1149, nx1151, nx1153, 
         nx1155, nx1157, nx1159, nx1161, nx1163, nx1165, nx1167, nx1169, nx1171, 
         nx1173, nx1175, nx1177, nx1179, nx1181, nx1183, nx1185, nx1187, nx1189, 
         nx1191, nx1193, nx1195, nx1197, nx1542, nx1544;



    OAI3R2 ix1259 (.X (l), .A1 (nx1248), .A2 (a[0]), .A3 (nx1195), .B (nx1197)
           ) ;
    OAI3R0 ix1249 (.X (nx1248), .A1 (nx1218), .A2 (nx1191), .A3 (b[1]), .B (
           nx1193)) ;
    OAI3R0 ix1219 (.X (nx1218), .A1 (nx1208), .A2 (a[2]), .A3 (nx1187), .B (
           nx1189)) ;
    OAI3R0 ix1209 (.X (nx1208), .A1 (nx1178), .A2 (nx1183), .A3 (b[3]), .B (
           nx1185)) ;
    OAI3R0 ix1179 (.X (nx1178), .A1 (nx1168), .A2 (a[4]), .A3 (nx1179), .B (
           nx1181)) ;
    OAI3R0 ix1169 (.X (nx1168), .A1 (nx1138), .A2 (nx1175), .A3 (b[5]), .B (
           nx1177)) ;
    OAI3R0 ix1139 (.X (nx1138), .A1 (nx1128), .A2 (a[6]), .A3 (nx1171), .B (
           nx1173)) ;
    OAI3R0 ix1129 (.X (nx1128), .A1 (nx1098), .A2 (nx1167), .A3 (b[7]), .B (
           nx1169)) ;
    OAI3R0 ix1099 (.X (nx1098), .A1 (nx1088), .A2 (a[8]), .A3 (nx1163), .B (
           nx1165)) ;
    OAI3R0 ix1089 (.X (nx1088), .A1 (nx1058), .A2 (nx1159), .A3 (b[9]), .B (
           nx1161)) ;
    OAI3R0 ix1059 (.X (nx1058), .A1 (nx1048), .A2 (a[10]), .A3 (nx1155), .B (
           nx1157)) ;
    OAI3R0 ix1049 (.X (nx1048), .A1 (nx1018), .A2 (nx1151), .A3 (b[11]), .B (
           nx1153)) ;
    OAI3R0 ix1019 (.X (nx1018), .A1 (nx1008), .A2 (a[12]), .A3 (nx1147), .B (
           nx1149)) ;
    OAI3R0 ix1009 (.X (nx1008), .A1 (nx978), .A2 (nx1143), .A3 (b[13]), .B (
           nx1145)) ;
    OAI3R0 ix979 (.X (nx978), .A1 (nx968), .A2 (a[14]), .A3 (nx1139), .B (nx1141
           )) ;
    OAI3R0 ix969 (.X (nx968), .A1 (nx938), .A2 (nx1135), .A3 (b[15]), .B (nx1137
           )) ;
    OAI3R0 ix939 (.X (nx938), .A1 (nx928), .A2 (a[16]), .A3 (nx1131), .B (nx1133
           )) ;
    OAI3R0 ix929 (.X (nx928), .A1 (nx898), .A2 (nx1127), .A3 (b[17]), .B (nx1129
           )) ;
    OAI3R0 ix899 (.X (nx898), .A1 (nx888), .A2 (a[18]), .A3 (nx1123), .B (nx1125
           )) ;
    OAI3R0 ix889 (.X (nx888), .A1 (nx858), .A2 (nx1119), .A3 (b[19]), .B (nx1121
           )) ;
    OAI3R0 ix859 (.X (nx858), .A1 (nx848), .A2 (a[20]), .A3 (nx1115), .B (nx1117
           )) ;
    OAI3R0 ix849 (.X (nx848), .A1 (nx818), .A2 (nx1111), .A3 (b[21]), .B (nx1113
           )) ;
    OAI3R0 ix819 (.X (nx818), .A1 (nx808), .A2 (a[22]), .A3 (nx1107), .B (nx1109
           )) ;
    OAI3R0 ix809 (.X (nx808), .A1 (nx778), .A2 (nx1103), .A3 (b[23]), .B (nx1105
           )) ;
    OAI3R0 ix779 (.X (nx778), .A1 (nx768), .A2 (a[24]), .A3 (nx1099), .B (nx1101
           )) ;
    OAI3R0 ix769 (.X (nx768), .A1 (nx738), .A2 (nx1095), .A3 (b[25]), .B (nx1097
           )) ;
    OAI3R0 ix739 (.X (nx738), .A1 (nx728), .A2 (a[26]), .A3 (nx1091), .B (nx1093
           )) ;
    OAI3R0 ix729 (.X (nx728), .A1 (nx698), .A2 (nx1087), .A3 (b[27]), .B (nx1089
           )) ;
    OAI3R0 ix699 (.X (nx698), .A1 (nx688), .A2 (a[28]), .A3 (nx1083), .B (nx1085
           )) ;
    OAI3R0 ix689 (.X (nx688), .A1 (nx658), .A2 (nx1079), .A3 (b[29]), .B (nx1081
           )) ;
    OAI3R0 ix659 (.X (nx658), .A1 (nx648), .A2 (a[30]), .A3 (nx1075), .B (nx1077
           )) ;
    OAI3R0 ix649 (.X (nx648), .A1 (nx618), .A2 (nx1071), .A3 (b[31]), .B (nx1073
           )) ;
    OAI3R0 ix619 (.X (nx618), .A1 (nx608), .A2 (a[32]), .A3 (nx1067), .B (nx1069
           )) ;
    OAI3R0 ix609 (.X (nx608), .A1 (nx578), .A2 (nx1063), .A3 (b[33]), .B (nx1065
           )) ;
    OAI3R0 ix579 (.X (nx578), .A1 (nx568), .A2 (a[34]), .A3 (nx1059), .B (nx1061
           )) ;
    OAI3R0 ix569 (.X (nx568), .A1 (nx538), .A2 (nx1055), .A3 (b[35]), .B (nx1057
           )) ;
    OAI3R0 ix539 (.X (nx538), .A1 (nx528), .A2 (a[36]), .A3 (nx1051), .B (nx1053
           )) ;
    OAI3R0 ix529 (.X (nx528), .A1 (nx498), .A2 (nx1047), .A3 (b[37]), .B (nx1049
           )) ;
    OAI3R0 ix499 (.X (nx498), .A1 (nx488), .A2 (a[38]), .A3 (nx1043), .B (nx1045
           )) ;
    OAI3R0 ix489 (.X (nx488), .A1 (nx458), .A2 (nx1039), .A3 (b[39]), .B (nx1041
           )) ;
    OAI3R0 ix459 (.X (nx458), .A1 (nx448), .A2 (a[40]), .A3 (nx1035), .B (nx1037
           )) ;
    OAI3R0 ix449 (.X (nx448), .A1 (nx418), .A2 (nx1031), .A3 (b[41]), .B (nx1033
           )) ;
    OAI3R0 ix419 (.X (nx418), .A1 (nx408), .A2 (a[42]), .A3 (nx1027), .B (nx1029
           )) ;
    OAI3R0 ix409 (.X (nx408), .A1 (nx378), .A2 (nx1023), .A3 (b[43]), .B (nx1025
           )) ;
    OAI3R0 ix379 (.X (nx378), .A1 (nx368), .A2 (a[44]), .A3 (nx1019), .B (nx1021
           )) ;
    OAI3R0 ix369 (.X (nx368), .A1 (nx338), .A2 (nx1015), .A3 (b[45]), .B (nx1017
           )) ;
    OAI3R0 ix339 (.X (nx338), .A1 (nx328), .A2 (a[46]), .A3 (nx1011), .B (nx1013
           )) ;
    OAI3R0 ix329 (.X (nx328), .A1 (nx298), .A2 (nx1007), .A3 (b[47]), .B (nx1009
           )) ;
    OAI3R0 ix299 (.X (nx298), .A1 (nx288), .A2 (a[48]), .A3 (nx1003), .B (nx1005
           )) ;
    OAI3R0 ix289 (.X (nx288), .A1 (nx258), .A2 (nx999), .A3 (b[49]), .B (nx1001)
           ) ;
    OAI3R0 ix259 (.X (nx258), .A1 (nx248), .A2 (a[50]), .A3 (nx995), .B (nx997)
           ) ;
    OAI3R0 ix249 (.X (nx248), .A1 (nx218), .A2 (nx991), .A3 (b[51]), .B (nx993)
           ) ;
    OAI3R0 ix219 (.X (nx218), .A1 (nx208), .A2 (a[52]), .A3 (nx987), .B (nx989)
           ) ;
    OAI3R0 ix209 (.X (nx208), .A1 (nx178), .A2 (nx983), .A3 (b[53]), .B (nx985)
           ) ;
    OAI3R0 ix179 (.X (nx178), .A1 (nx168), .A2 (a[54]), .A3 (nx979), .B (nx981)
           ) ;
    OAI3R0 ix169 (.X (nx168), .A1 (nx138), .A2 (nx975), .A3 (b[55]), .B (nx977)
           ) ;
    OAI3R0 ix139 (.X (nx138), .A1 (nx128), .A2 (a[56]), .A3 (nx971), .B (nx973)
           ) ;
    OAI3R0 ix129 (.X (nx128), .A1 (nx98), .A2 (nx967), .A3 (b[57]), .B (nx969)
           ) ;
    OAI3R0 ix99 (.X (nx98), .A1 (nx88), .A2 (a[58]), .A3 (nx963), .B (nx965)) ;
    OAI3R0 ix89 (.X (nx88), .A1 (nx58), .A2 (nx959), .A3 (b[59]), .B (nx961)) ;
    OAI3R0 ix59 (.X (nx58), .A1 (nx48), .A2 (a[60]), .A3 (nx955), .B (nx957)) ;
    OAI3R0 ix49 (.X (nx48), .A1 (nx28), .A2 (nx947), .A3 (b[61]), .B (nx949)) ;
    OAI1A0 ix29 (.X (nx28), .A1 (a[63]), .A2 (nx939), .B (nx941)) ;
    IV1N0 ix940 (.X (nx939), .A (b[63])) ;
    OAI3N0 ix942 (.X (nx941), .A1 (nx943), .A2 (b[63]), .B1 (nx945), .B2 (b[62])
           ) ;
    IV1N0 ix944 (.X (nx943), .A (a[63])) ;
    IV1N0 ix946 (.X (nx945), .A (a[62])) ;
    IV1N0 ix948 (.X (nx947), .A (a[61])) ;
    OAI3N0 ix952 (.X (nx951), .A1 (nx939), .A2 (a[63]), .B1 (a[62]), .B2 (nx953)
           ) ;
    IV1N0 ix954 (.X (nx953), .A (b[62])) ;
    IV1N0 ix956 (.X (nx955), .A (b[60])) ;
    AO3I0 ix958 (.X (nx957), .A1 (nx949), .A2 (nx947), .A3 (b[61]), .B (nx28)) ;
    IV1N0 ix960 (.X (nx959), .A (a[59])) ;
    AO3I0 ix962 (.X (nx961), .A1 (nx957), .A2 (a[60]), .A3 (nx955), .B (nx48)) ;
    IV1N0 ix964 (.X (nx963), .A (b[58])) ;
    AO3I0 ix966 (.X (nx965), .A1 (nx961), .A2 (nx959), .A3 (b[59]), .B (nx58)) ;
    IV1N0 ix968 (.X (nx967), .A (a[57])) ;
    AO3I0 ix970 (.X (nx969), .A1 (nx965), .A2 (a[58]), .A3 (nx963), .B (nx88)) ;
    IV1N0 ix972 (.X (nx971), .A (b[56])) ;
    AO3I0 ix974 (.X (nx973), .A1 (nx969), .A2 (nx967), .A3 (b[57]), .B (nx98)) ;
    IV1N0 ix976 (.X (nx975), .A (a[55])) ;
    AO3I0 ix978 (.X (nx977), .A1 (nx973), .A2 (a[56]), .A3 (nx971), .B (nx128)
          ) ;
    IV1N0 ix980 (.X (nx979), .A (b[54])) ;
    AO3I0 ix982 (.X (nx981), .A1 (nx977), .A2 (nx975), .A3 (b[55]), .B (nx138)
          ) ;
    IV1N0 ix984 (.X (nx983), .A (a[53])) ;
    AO3I0 ix986 (.X (nx985), .A1 (nx981), .A2 (a[54]), .A3 (nx979), .B (nx168)
          ) ;
    IV1N0 ix988 (.X (nx987), .A (b[52])) ;
    AO3I0 ix990 (.X (nx989), .A1 (nx985), .A2 (nx983), .A3 (b[53]), .B (nx178)
          ) ;
    IV1N0 ix992 (.X (nx991), .A (a[51])) ;
    AO3I0 ix994 (.X (nx993), .A1 (nx989), .A2 (a[52]), .A3 (nx987), .B (nx208)
          ) ;
    IV1N0 ix996 (.X (nx995), .A (b[50])) ;
    AO3I0 ix998 (.X (nx997), .A1 (nx993), .A2 (nx991), .A3 (b[51]), .B (nx218)
          ) ;
    IV1N0 ix1000 (.X (nx999), .A (a[49])) ;
    AO3I0 ix1002 (.X (nx1001), .A1 (nx997), .A2 (a[50]), .A3 (nx995), .B (nx248)
          ) ;
    IV1N0 ix1004 (.X (nx1003), .A (b[48])) ;
    AO3I0 ix1006 (.X (nx1005), .A1 (nx1001), .A2 (nx999), .A3 (b[49]), .B (nx258
          )) ;
    IV1N0 ix1008 (.X (nx1007), .A (a[47])) ;
    AO3I0 ix1010 (.X (nx1009), .A1 (nx1005), .A2 (a[48]), .A3 (nx1003), .B (
          nx288)) ;
    IV1N0 ix1012 (.X (nx1011), .A (b[46])) ;
    AO3I0 ix1014 (.X (nx1013), .A1 (nx1009), .A2 (nx1007), .A3 (b[47]), .B (
          nx298)) ;
    IV1N0 ix1016 (.X (nx1015), .A (a[45])) ;
    AO3I0 ix1018 (.X (nx1017), .A1 (nx1013), .A2 (a[46]), .A3 (nx1011), .B (
          nx328)) ;
    IV1N0 ix1020 (.X (nx1019), .A (b[44])) ;
    AO3I0 ix1022 (.X (nx1021), .A1 (nx1017), .A2 (nx1015), .A3 (b[45]), .B (
          nx338)) ;
    IV1N0 ix1024 (.X (nx1023), .A (a[43])) ;
    AO3I0 ix1026 (.X (nx1025), .A1 (nx1021), .A2 (a[44]), .A3 (nx1019), .B (
          nx368)) ;
    IV1N0 ix1028 (.X (nx1027), .A (b[42])) ;
    AO3I0 ix1030 (.X (nx1029), .A1 (nx1025), .A2 (nx1023), .A3 (b[43]), .B (
          nx378)) ;
    IV1N0 ix1032 (.X (nx1031), .A (a[41])) ;
    AO3I0 ix1034 (.X (nx1033), .A1 (nx1029), .A2 (a[42]), .A3 (nx1027), .B (
          nx408)) ;
    IV1N0 ix1036 (.X (nx1035), .A (b[40])) ;
    AO3I0 ix1038 (.X (nx1037), .A1 (nx1033), .A2 (nx1031), .A3 (b[41]), .B (
          nx418)) ;
    IV1N0 ix1040 (.X (nx1039), .A (a[39])) ;
    AO3I0 ix1042 (.X (nx1041), .A1 (nx1037), .A2 (a[40]), .A3 (nx1035), .B (
          nx448)) ;
    IV1N0 ix1044 (.X (nx1043), .A (b[38])) ;
    AO3I0 ix1046 (.X (nx1045), .A1 (nx1041), .A2 (nx1039), .A3 (b[39]), .B (
          nx458)) ;
    IV1N0 ix1048 (.X (nx1047), .A (a[37])) ;
    AO3I0 ix1050 (.X (nx1049), .A1 (nx1045), .A2 (a[38]), .A3 (nx1043), .B (
          nx488)) ;
    IV1N0 ix1052 (.X (nx1051), .A (b[36])) ;
    AO3I0 ix1054 (.X (nx1053), .A1 (nx1049), .A2 (nx1047), .A3 (b[37]), .B (
          nx498)) ;
    IV1N0 ix1056 (.X (nx1055), .A (a[35])) ;
    AO3I0 ix1058 (.X (nx1057), .A1 (nx1053), .A2 (a[36]), .A3 (nx1051), .B (
          nx528)) ;
    IV1N0 ix1060 (.X (nx1059), .A (b[34])) ;
    AO3I0 ix1062 (.X (nx1061), .A1 (nx1057), .A2 (nx1055), .A3 (b[35]), .B (
          nx538)) ;
    IV1N0 ix1064 (.X (nx1063), .A (a[33])) ;
    AO3I0 ix1066 (.X (nx1065), .A1 (nx1061), .A2 (a[34]), .A3 (nx1059), .B (
          nx568)) ;
    IV1N0 ix1068 (.X (nx1067), .A (b[32])) ;
    AO3I0 ix1070 (.X (nx1069), .A1 (nx1065), .A2 (nx1063), .A3 (b[33]), .B (
          nx578)) ;
    IV1N0 ix1072 (.X (nx1071), .A (a[31])) ;
    AO3I0 ix1074 (.X (nx1073), .A1 (nx1069), .A2 (a[32]), .A3 (nx1067), .B (
          nx608)) ;
    IV1N0 ix1076 (.X (nx1075), .A (b[30])) ;
    AO3I0 ix1078 (.X (nx1077), .A1 (nx1073), .A2 (nx1071), .A3 (b[31]), .B (
          nx618)) ;
    IV1N0 ix1080 (.X (nx1079), .A (a[29])) ;
    AO3I0 ix1082 (.X (nx1081), .A1 (nx1077), .A2 (a[30]), .A3 (nx1075), .B (
          nx648)) ;
    IV1N0 ix1084 (.X (nx1083), .A (b[28])) ;
    AO3I0 ix1086 (.X (nx1085), .A1 (nx1081), .A2 (nx1079), .A3 (b[29]), .B (
          nx658)) ;
    IV1N0 ix1088 (.X (nx1087), .A (a[27])) ;
    AO3I0 ix1090 (.X (nx1089), .A1 (nx1085), .A2 (a[28]), .A3 (nx1083), .B (
          nx688)) ;
    IV1N0 ix1092 (.X (nx1091), .A (b[26])) ;
    AO3I0 ix1094 (.X (nx1093), .A1 (nx1089), .A2 (nx1087), .A3 (b[27]), .B (
          nx698)) ;
    IV1N0 ix1096 (.X (nx1095), .A (a[25])) ;
    AO3I0 ix1098 (.X (nx1097), .A1 (nx1093), .A2 (a[26]), .A3 (nx1091), .B (
          nx728)) ;
    IV1N0 ix1100 (.X (nx1099), .A (b[24])) ;
    AO3I0 ix1102 (.X (nx1101), .A1 (nx1097), .A2 (nx1095), .A3 (b[25]), .B (
          nx738)) ;
    IV1N0 ix1104 (.X (nx1103), .A (a[23])) ;
    AO3I0 ix1106 (.X (nx1105), .A1 (nx1101), .A2 (a[24]), .A3 (nx1099), .B (
          nx768)) ;
    IV1N0 ix1108 (.X (nx1107), .A (b[22])) ;
    AO3I0 ix1110 (.X (nx1109), .A1 (nx1105), .A2 (nx1103), .A3 (b[23]), .B (
          nx778)) ;
    IV1N0 ix1112 (.X (nx1111), .A (a[21])) ;
    AO3I0 ix1114 (.X (nx1113), .A1 (nx1109), .A2 (a[22]), .A3 (nx1107), .B (
          nx808)) ;
    IV1N0 ix1116 (.X (nx1115), .A (b[20])) ;
    AO3I0 ix1118 (.X (nx1117), .A1 (nx1113), .A2 (nx1111), .A3 (b[21]), .B (
          nx818)) ;
    IV1N0 ix1120 (.X (nx1119), .A (a[19])) ;
    AO3I0 ix1122 (.X (nx1121), .A1 (nx1117), .A2 (a[20]), .A3 (nx1115), .B (
          nx848)) ;
    IV1N0 ix1124 (.X (nx1123), .A (b[18])) ;
    AO3I0 ix1126 (.X (nx1125), .A1 (nx1121), .A2 (nx1119), .A3 (b[19]), .B (
          nx858)) ;
    IV1N0 ix1128 (.X (nx1127), .A (a[17])) ;
    AO3I0 ix1130 (.X (nx1129), .A1 (nx1125), .A2 (a[18]), .A3 (nx1123), .B (
          nx888)) ;
    IV1N0 ix1132 (.X (nx1131), .A (b[16])) ;
    AO3I0 ix1134 (.X (nx1133), .A1 (nx1129), .A2 (nx1127), .A3 (b[17]), .B (
          nx898)) ;
    IV1N0 ix1136 (.X (nx1135), .A (a[15])) ;
    AO3I0 ix1138 (.X (nx1137), .A1 (nx1133), .A2 (a[16]), .A3 (nx1131), .B (
          nx928)) ;
    IV1N0 ix1140 (.X (nx1139), .A (b[14])) ;
    AO3I0 ix1142 (.X (nx1141), .A1 (nx1137), .A2 (nx1135), .A3 (b[15]), .B (
          nx938)) ;
    IV1N0 ix1144 (.X (nx1143), .A (a[13])) ;
    AO3I0 ix1146 (.X (nx1145), .A1 (nx1141), .A2 (a[14]), .A3 (nx1139), .B (
          nx968)) ;
    IV1N0 ix1148 (.X (nx1147), .A (b[12])) ;
    AO3I0 ix1150 (.X (nx1149), .A1 (nx1145), .A2 (nx1143), .A3 (b[13]), .B (
          nx978)) ;
    IV1N0 ix1152 (.X (nx1151), .A (a[11])) ;
    AO3I0 ix1154 (.X (nx1153), .A1 (nx1149), .A2 (a[12]), .A3 (nx1147), .B (
          nx1008)) ;
    IV1N0 ix1156 (.X (nx1155), .A (b[10])) ;
    AO3I0 ix1158 (.X (nx1157), .A1 (nx1153), .A2 (nx1151), .A3 (b[11]), .B (
          nx1018)) ;
    IV1N0 ix1160 (.X (nx1159), .A (a[9])) ;
    AO3I0 ix1162 (.X (nx1161), .A1 (nx1157), .A2 (a[10]), .A3 (nx1155), .B (
          nx1048)) ;
    IV1N0 ix1164 (.X (nx1163), .A (b[8])) ;
    AO3I0 ix1166 (.X (nx1165), .A1 (nx1161), .A2 (nx1159), .A3 (b[9]), .B (
          nx1058)) ;
    IV1N0 ix1168 (.X (nx1167), .A (a[7])) ;
    AO3I0 ix1170 (.X (nx1169), .A1 (nx1165), .A2 (a[8]), .A3 (nx1163), .B (
          nx1088)) ;
    IV1N0 ix1172 (.X (nx1171), .A (b[6])) ;
    AO3I0 ix1174 (.X (nx1173), .A1 (nx1169), .A2 (nx1167), .A3 (b[7]), .B (
          nx1098)) ;
    IV1N0 ix1176 (.X (nx1175), .A (a[5])) ;
    AO3I0 ix1178 (.X (nx1177), .A1 (nx1173), .A2 (a[6]), .A3 (nx1171), .B (
          nx1128)) ;
    IV1N0 ix1180 (.X (nx1179), .A (b[4])) ;
    AO3I0 ix1182 (.X (nx1181), .A1 (nx1177), .A2 (nx1175), .A3 (b[5]), .B (
          nx1138)) ;
    IV1N0 ix1184 (.X (nx1183), .A (a[3])) ;
    AO3I0 ix1186 (.X (nx1185), .A1 (nx1181), .A2 (a[4]), .A3 (nx1179), .B (
          nx1168)) ;
    IV1N0 ix1188 (.X (nx1187), .A (b[2])) ;
    AO3I0 ix1190 (.X (nx1189), .A1 (nx1185), .A2 (nx1183), .A3 (b[3]), .B (
          nx1178)) ;
    IV1N0 ix1192 (.X (nx1191), .A (a[1])) ;
    AO3I0 ix1194 (.X (nx1193), .A1 (nx1189), .A2 (a[2]), .A3 (nx1187), .B (
          nx1208)) ;
    IV1N0 ix1196 (.X (nx1195), .A (b[0])) ;
    AO3I0 ix1198 (.X (nx1197), .A1 (nx1193), .A2 (nx1191), .A3 (b[1]), .B (
          nx1218)) ;
    OAI3R0 ix1269 (.X (g), .A1 (nx1238), .A2 (nx1542), .A3 (b[0]), .B (nx1544)
           ) ;
    IV1N0 ix1543 (.X (nx1542), .A (a[0])) ;
    IV1N0 ix1545 (.X (nx1544), .A (nx1248)) ;
    IV1N0 ix1239 (.X (nx1238), .A (nx1197)) ;
    OA1R0 ix15 (.X (nx949), .A1 (nx943), .A2 (b[63]), .B (nx951)) ;
endmodule


module OA1R0 ( X, A1, A2, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input B ;

    wire nx0, nx2;



    and (nx0, A2, B) ;
    and (nx2, A1, B) ;
    or (X, nx0, nx2) ;
endmodule


module AO3I0 ( X, A1, A2, A3, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input A3 ;
    input B ;

    wire NOT_A3, NOT_B, nx4, NOT_A2, nx8, nx10, NOT_A1, nx14;



    assign NOT_A3 = ~A3 ;
    assign NOT_B = ~B ;
    and (nx4, NOT_A3, NOT_B) ;
    assign NOT_A2 = ~A2 ;
    and (nx8, NOT_A2, NOT_B) ;
    or (nx10, nx4, nx8) ;
    assign NOT_A1 = ~A1 ;
    and (nx14, NOT_A1, NOT_B) ;
    or (X, nx10, nx14) ;
endmodule


module OAI3N0 ( X, A1, A2, B1, B2 ) ;

    output X ;
    input A1 ;
    input A2 ;
    input B1 ;
    input B2 ;

    wire NOT_A1, NOT_A2, nx4, NOT_B2, nx8, NOT_B1;



    assign NOT_A1 = ~A1 ;
    assign NOT_A2 = ~A2 ;
    and (nx4, NOT_A1, NOT_A2) ;
    assign NOT_B2 = ~B2 ;
    or (nx8, nx4, NOT_B2) ;
    assign NOT_B1 = ~B1 ;
    or (X, nx8, NOT_B1) ;
endmodule


module IV1N0 ( X, A ) ;

    output X ;
    input A ;




    assign X = ~A ;
endmodule


module OAI1A0 ( X, A1, A2, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input B ;

    wire NOT_A1, NOT_A2, nx4, NOT_B;



    assign NOT_A1 = ~A1 ;
    assign NOT_A2 = ~A2 ;
    and (nx4, NOT_A1, NOT_A2) ;
    assign NOT_B = ~B ;
    or (X, nx4, NOT_B) ;
endmodule


module OAI3R0 ( X, A1, A2, A3, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input A3 ;
    input B ;

    wire NOT_A1, NOT_A2, nx4, NOT_A3, nx8, NOT_B;



    assign NOT_A1 = ~A1 ;
    assign NOT_A2 = ~A2 ;
    and (nx4, NOT_A1, NOT_A2) ;
    assign NOT_A3 = ~A3 ;
    and (nx8, nx4, NOT_A3) ;
    assign NOT_B = ~B ;
    or (X, nx8, NOT_B) ;
endmodule


module OAI3R2 ( X, A1, A2, A3, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input A3 ;
    input B ;

    wire NOT_A1, NOT_A2, nx4, NOT_A3, nx8, NOT_B;



    assign NOT_A1 = ~A1 ;
    assign NOT_A2 = ~A2 ;
    and (nx4, NOT_A1, NOT_A2) ;
    assign NOT_A3 = ~A3 ;
    and (nx8, nx4, NOT_A3) ;
    assign NOT_B = ~B ;
    or (X, nx8, NOT_B) ;
endmodule

