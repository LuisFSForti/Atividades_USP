* C:\Users\luis\Documents\Facul\Atividades_USP\Circuitos\EX3\14592348.sch

* Schematics Version 9.1 - Web Update 1
* Thu Jun 27 17:22:06 2024



** Analysis setup **
.tran 10us 1


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "14592348.net"
.INC "14592348.als"


.probe


.END
