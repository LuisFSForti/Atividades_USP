//
// Verilog description for cell ordenador, 
// 06/12/24 10:25:34
//
// LeonardoSpectrum Level 3, 2020a.2 
//


module ordenador ( y8, y7, y6, y5, y4, y3, y2, y1, x8, x7, x6, x5, x4, x3, x2, 
                   x1 ) ;

    output [31:0]y8 ;
    output [31:0]y7 ;
    output [31:0]y6 ;
    output [31:0]y5 ;
    output [31:0]y4 ;
    output [31:0]y3 ;
    output [31:0]y2 ;
    output [31:0]y1 ;
    input [31:0]x8 ;
    input [31:0]x7 ;
    input [31:0]x6 ;
    input [31:0]x5 ;
    input [31:0]x4 ;
    input [31:0]x3 ;
    input [31:0]x2 ;
    input [31:0]x1 ;

    wire linha7_7__31, linha7_7__30, linha7_7__29, linha7_7__28, linha7_7__27, 
         linha7_7__26, linha7_7__25, linha7_7__24, linha7_7__23, linha7_7__22, 
         linha7_7__21, linha7_7__20, linha7_7__19, linha7_7__18, linha7_7__17, 
         linha7_7__16, linha7_7__15, linha7_7__14, linha7_7__13, linha7_7__12, 
         linha7_7__11, linha7_7__10, linha7_7__9, linha7_7__8, linha7_7__7, 
         linha7_7__6, linha7_7__5, linha7_7__4, linha7_7__3, linha7_7__2, 
         linha7_7__1, linha7_7__0, linha7_6__31, linha7_6__30, linha7_6__29, 
         linha7_6__28, linha7_6__27, linha7_6__26, linha7_6__25, linha7_6__24, 
         linha7_6__23, linha7_6__22, linha7_6__21, linha7_6__20, linha7_6__19, 
         linha7_6__18, linha7_6__17, linha7_6__16, linha7_6__15, linha7_6__14, 
         linha7_6__13, linha7_6__12, linha7_6__11, linha7_6__10, linha7_6__9, 
         linha7_6__8, linha7_6__7, linha7_6__6, linha7_6__5, linha7_6__4, 
         linha7_6__3, linha7_6__2, linha7_6__1, linha7_6__0, linha7_5__31, 
         linha7_5__30, linha7_5__29, linha7_5__28, linha7_5__27, linha7_5__26, 
         linha7_5__25, linha7_5__24, linha7_5__23, linha7_5__22, linha7_5__21, 
         linha7_5__20, linha7_5__19, linha7_5__18, linha7_5__17, linha7_5__16, 
         linha7_5__15, linha7_5__14, linha7_5__13, linha7_5__12, linha7_5__11, 
         linha7_5__10, linha7_5__9, linha7_5__8, linha7_5__7, linha7_5__6, 
         linha7_5__5, linha7_5__4, linha7_5__3, linha7_5__2, linha7_5__1, 
         linha7_5__0, linha7_4__31, linha7_4__30, linha7_4__29, linha7_4__28, 
         linha7_4__27, linha7_4__26, linha7_4__25, linha7_4__24, linha7_4__23, 
         linha7_4__22, linha7_4__21, linha7_4__20, linha7_4__19, linha7_4__18, 
         linha7_4__17, linha7_4__16, linha7_4__15, linha7_4__14, linha7_4__13, 
         linha7_4__12, linha7_4__11, linha7_4__10, linha7_4__9, linha7_4__8, 
         linha7_4__7, linha7_4__6, linha7_4__5, linha7_4__4, linha7_4__3, 
         linha7_4__2, linha7_4__1, linha7_4__0, linha7_3__31, linha7_3__30, 
         linha7_3__29, linha7_3__28, linha7_3__27, linha7_3__26, linha7_3__25, 
         linha7_3__24, linha7_3__23, linha7_3__22, linha7_3__21, linha7_3__20, 
         linha7_3__19, linha7_3__18, linha7_3__17, linha7_3__16, linha7_3__15, 
         linha7_3__14, linha7_3__13, linha7_3__12, linha7_3__11, linha7_3__10, 
         linha7_3__9, linha7_3__8, linha7_3__7, linha7_3__6, linha7_3__5, 
         linha7_3__4, linha7_3__3, linha7_3__2, linha7_3__1, linha7_3__0, 
         linha7_2__31, linha7_2__30, linha7_2__29, linha7_2__28, linha7_2__27, 
         linha7_2__26, linha7_2__25, linha7_2__24, linha7_2__23, linha7_2__22, 
         linha7_2__21, linha7_2__20, linha7_2__19, linha7_2__18, linha7_2__17, 
         linha7_2__16, linha7_2__15, linha7_2__14, linha7_2__13, linha7_2__12, 
         linha7_2__11, linha7_2__10, linha7_2__9, linha7_2__8, linha7_2__7, 
         linha7_2__6, linha7_2__5, linha7_2__4, linha7_2__3, linha7_2__2, 
         linha7_2__1, linha7_2__0, linha7_1__31, linha7_1__30, linha7_1__29, 
         linha7_1__28, linha7_1__27, linha7_1__26, linha7_1__25, linha7_1__24, 
         linha7_1__23, linha7_1__22, linha7_1__21, linha7_1__20, linha7_1__19, 
         linha7_1__18, linha7_1__17, linha7_1__16, linha7_1__15, linha7_1__14, 
         linha7_1__13, linha7_1__12, linha7_1__11, linha7_1__10, linha7_1__9, 
         linha7_1__8, linha7_1__7, linha7_1__6, linha7_1__5, linha7_1__4, 
         linha7_1__3, linha7_1__2, linha7_1__1, linha7_1__0, linha6_7__31, 
         linha6_7__30, linha6_7__29, linha6_7__28, linha6_7__27, linha6_7__26, 
         linha6_7__25, linha6_7__24, linha6_7__23, linha6_7__22, linha6_7__21, 
         linha6_7__20, linha6_7__19, linha6_7__18, linha6_7__17, linha6_7__16, 
         linha6_7__15, linha6_7__14, linha6_7__13, linha6_7__12, linha6_7__11, 
         linha6_7__10, linha6_7__9, linha6_7__8, linha6_7__7, linha6_7__6, 
         linha6_7__5, linha6_7__4, linha6_7__3, linha6_7__2, linha6_7__1, 
         linha6_7__0, linha6_6__31, linha6_6__30, linha6_6__29, linha6_6__28, 
         linha6_6__27, linha6_6__26, linha6_6__25, linha6_6__24, linha6_6__23, 
         linha6_6__22, linha6_6__21, linha6_6__20, linha6_6__19, linha6_6__18, 
         linha6_6__17, linha6_6__16, linha6_6__15, linha6_6__14, linha6_6__13, 
         linha6_6__12, linha6_6__11, linha6_6__10, linha6_6__9, linha6_6__8, 
         linha6_6__7, linha6_6__6, linha6_6__5, linha6_6__4, linha6_6__3, 
         linha6_6__2, linha6_6__1, linha6_6__0, linha6_5__31, linha6_5__30, 
         linha6_5__29, linha6_5__28, linha6_5__27, linha6_5__26, linha6_5__25, 
         linha6_5__24, linha6_5__23, linha6_5__22, linha6_5__21, linha6_5__20, 
         linha6_5__19, linha6_5__18, linha6_5__17, linha6_5__16, linha6_5__15, 
         linha6_5__14, linha6_5__13, linha6_5__12, linha6_5__11, linha6_5__10, 
         linha6_5__9, linha6_5__8, linha6_5__7, linha6_5__6, linha6_5__5, 
         linha6_5__4, linha6_5__3, linha6_5__2, linha6_5__1, linha6_5__0, 
         linha6_4__31, linha6_4__30, linha6_4__29, linha6_4__28, linha6_4__27, 
         linha6_4__26, linha6_4__25, linha6_4__24, linha6_4__23, linha6_4__22, 
         linha6_4__21, linha6_4__20, linha6_4__19, linha6_4__18, linha6_4__17, 
         linha6_4__16, linha6_4__15, linha6_4__14, linha6_4__13, linha6_4__12, 
         linha6_4__11, linha6_4__10, linha6_4__9, linha6_4__8, linha6_4__7, 
         linha6_4__6, linha6_4__5, linha6_4__4, linha6_4__3, linha6_4__2, 
         linha6_4__1, linha6_4__0, linha6_3__31, linha6_3__30, linha6_3__29, 
         linha6_3__28, linha6_3__27, linha6_3__26, linha6_3__25, linha6_3__24, 
         linha6_3__23, linha6_3__22, linha6_3__21, linha6_3__20, linha6_3__19, 
         linha6_3__18, linha6_3__17, linha6_3__16, linha6_3__15, linha6_3__14, 
         linha6_3__13, linha6_3__12, linha6_3__11, linha6_3__10, linha6_3__9, 
         linha6_3__8, linha6_3__7, linha6_3__6, linha6_3__5, linha6_3__4, 
         linha6_3__3, linha6_3__2, linha6_3__1, linha6_3__0, linha6_2__31, 
         linha6_2__30, linha6_2__29, linha6_2__28, linha6_2__27, linha6_2__26, 
         linha6_2__25, linha6_2__24, linha6_2__23, linha6_2__22, linha6_2__21, 
         linha6_2__20, linha6_2__19, linha6_2__18, linha6_2__17, linha6_2__16, 
         linha6_2__15, linha6_2__14, linha6_2__13, linha6_2__12, linha6_2__11, 
         linha6_2__10, linha6_2__9, linha6_2__8, linha6_2__7, linha6_2__6, 
         linha6_2__5, linha6_2__4, linha6_2__3, linha6_2__2, linha6_2__1, 
         linha6_2__0, linha6_1__31, linha6_1__30, linha6_1__29, linha6_1__28, 
         linha6_1__27, linha6_1__26, linha6_1__25, linha6_1__24, linha6_1__23, 
         linha6_1__22, linha6_1__21, linha6_1__20, linha6_1__19, linha6_1__18, 
         linha6_1__17, linha6_1__16, linha6_1__15, linha6_1__14, linha6_1__13, 
         linha6_1__12, linha6_1__11, linha6_1__10, linha6_1__9, linha6_1__8, 
         linha6_1__7, linha6_1__6, linha6_1__5, linha6_1__4, linha6_1__3, 
         linha6_1__2, linha6_1__1, linha6_1__0, linha5_7__31, linha5_7__30, 
         linha5_7__29, linha5_7__28, linha5_7__27, linha5_7__26, linha5_7__25, 
         linha5_7__24, linha5_7__23, linha5_7__22, linha5_7__21, linha5_7__20, 
         linha5_7__19, linha5_7__18, linha5_7__17, linha5_7__16, linha5_7__15, 
         linha5_7__14, linha5_7__13, linha5_7__12, linha5_7__11, linha5_7__10, 
         linha5_7__9, linha5_7__8, linha5_7__7, linha5_7__6, linha5_7__5, 
         linha5_7__4, linha5_7__3, linha5_7__2, linha5_7__1, linha5_7__0, 
         linha5_6__31, linha5_6__30, linha5_6__29, linha5_6__28, linha5_6__27, 
         linha5_6__26, linha5_6__25, linha5_6__24, linha5_6__23, linha5_6__22, 
         linha5_6__21, linha5_6__20, linha5_6__19, linha5_6__18, linha5_6__17, 
         linha5_6__16, linha5_6__15, linha5_6__14, linha5_6__13, linha5_6__12, 
         linha5_6__11, linha5_6__10, linha5_6__9, linha5_6__8, linha5_6__7, 
         linha5_6__6, linha5_6__5, linha5_6__4, linha5_6__3, linha5_6__2, 
         linha5_6__1, linha5_6__0, linha5_5__31, linha5_5__30, linha5_5__29, 
         linha5_5__28, linha5_5__27, linha5_5__26, linha5_5__25, linha5_5__24, 
         linha5_5__23, linha5_5__22, linha5_5__21, linha5_5__20, linha5_5__19, 
         linha5_5__18, linha5_5__17, linha5_5__16, linha5_5__15, linha5_5__14, 
         linha5_5__13, linha5_5__12, linha5_5__11, linha5_5__10, linha5_5__9, 
         linha5_5__8, linha5_5__7, linha5_5__6, linha5_5__5, linha5_5__4, 
         linha5_5__3, linha5_5__2, linha5_5__1, linha5_5__0, linha5_4__31, 
         linha5_4__30, linha5_4__29, linha5_4__28, linha5_4__27, linha5_4__26, 
         linha5_4__25, linha5_4__24, linha5_4__23, linha5_4__22, linha5_4__21, 
         linha5_4__20, linha5_4__19, linha5_4__18, linha5_4__17, linha5_4__16, 
         linha5_4__15, linha5_4__14, linha5_4__13, linha5_4__12, linha5_4__11, 
         linha5_4__10, linha5_4__9, linha5_4__8, linha5_4__7, linha5_4__6, 
         linha5_4__5, linha5_4__4, linha5_4__3, linha5_4__2, linha5_4__1, 
         linha5_4__0, linha5_3__31, linha5_3__30, linha5_3__29, linha5_3__28, 
         linha5_3__27, linha5_3__26, linha5_3__25, linha5_3__24, linha5_3__23, 
         linha5_3__22, linha5_3__21, linha5_3__20, linha5_3__19, linha5_3__18, 
         linha5_3__17, linha5_3__16, linha5_3__15, linha5_3__14, linha5_3__13, 
         linha5_3__12, linha5_3__11, linha5_3__10, linha5_3__9, linha5_3__8, 
         linha5_3__7, linha5_3__6, linha5_3__5, linha5_3__4, linha5_3__3, 
         linha5_3__2, linha5_3__1, linha5_3__0, linha5_2__31, linha5_2__30, 
         linha5_2__29, linha5_2__28, linha5_2__27, linha5_2__26, linha5_2__25, 
         linha5_2__24, linha5_2__23, linha5_2__22, linha5_2__21, linha5_2__20, 
         linha5_2__19, linha5_2__18, linha5_2__17, linha5_2__16, linha5_2__15, 
         linha5_2__14, linha5_2__13, linha5_2__12, linha5_2__11, linha5_2__10, 
         linha5_2__9, linha5_2__8, linha5_2__7, linha5_2__6, linha5_2__5, 
         linha5_2__4, linha5_2__3, linha5_2__2, linha5_2__1, linha5_2__0, 
         linha5_1__31, linha5_1__30, linha5_1__29, linha5_1__28, linha5_1__27, 
         linha5_1__26, linha5_1__25, linha5_1__24, linha5_1__23, linha5_1__22, 
         linha5_1__21, linha5_1__20, linha5_1__19, linha5_1__18, linha5_1__17, 
         linha5_1__16, linha5_1__15, linha5_1__14, linha5_1__13, linha5_1__12, 
         linha5_1__11, linha5_1__10, linha5_1__9, linha5_1__8, linha5_1__7, 
         linha5_1__6, linha5_1__5, linha5_1__4, linha5_1__3, linha5_1__2, 
         linha5_1__1, linha5_1__0, linha4_7__31, linha4_7__30, linha4_7__29, 
         linha4_7__28, linha4_7__27, linha4_7__26, linha4_7__25, linha4_7__24, 
         linha4_7__23, linha4_7__22, linha4_7__21, linha4_7__20, linha4_7__19, 
         linha4_7__18, linha4_7__17, linha4_7__16, linha4_7__15, linha4_7__14, 
         linha4_7__13, linha4_7__12, linha4_7__11, linha4_7__10, linha4_7__9, 
         linha4_7__8, linha4_7__7, linha4_7__6, linha4_7__5, linha4_7__4, 
         linha4_7__3, linha4_7__2, linha4_7__1, linha4_7__0, linha4_6__31, 
         linha4_6__30, linha4_6__29, linha4_6__28, linha4_6__27, linha4_6__26, 
         linha4_6__25, linha4_6__24, linha4_6__23, linha4_6__22, linha4_6__21, 
         linha4_6__20, linha4_6__19, linha4_6__18, linha4_6__17, linha4_6__16, 
         linha4_6__15, linha4_6__14, linha4_6__13, linha4_6__12, linha4_6__11, 
         linha4_6__10, linha4_6__9, linha4_6__8, linha4_6__7, linha4_6__6, 
         linha4_6__5, linha4_6__4, linha4_6__3, linha4_6__2, linha4_6__1, 
         linha4_6__0, linha4_5__31, linha4_5__30, linha4_5__29, linha4_5__28, 
         linha4_5__27, linha4_5__26, linha4_5__25, linha4_5__24, linha4_5__23, 
         linha4_5__22, linha4_5__21, linha4_5__20, linha4_5__19, linha4_5__18, 
         linha4_5__17, linha4_5__16, linha4_5__15, linha4_5__14, linha4_5__13, 
         linha4_5__12, linha4_5__11, linha4_5__10, linha4_5__9, linha4_5__8, 
         linha4_5__7, linha4_5__6, linha4_5__5, linha4_5__4, linha4_5__3, 
         linha4_5__2, linha4_5__1, linha4_5__0, linha4_4__31, linha4_4__30, 
         linha4_4__29, linha4_4__28, linha4_4__27, linha4_4__26, linha4_4__25, 
         linha4_4__24, linha4_4__23, linha4_4__22, linha4_4__21, linha4_4__20, 
         linha4_4__19, linha4_4__18, linha4_4__17, linha4_4__16, linha4_4__15, 
         linha4_4__14, linha4_4__13, linha4_4__12, linha4_4__11, linha4_4__10, 
         linha4_4__9, linha4_4__8, linha4_4__7, linha4_4__6, linha4_4__5, 
         linha4_4__4, linha4_4__3, linha4_4__2, linha4_4__1, linha4_4__0, 
         linha4_3__31, linha4_3__30, linha4_3__29, linha4_3__28, linha4_3__27, 
         linha4_3__26, linha4_3__25, linha4_3__24, linha4_3__23, linha4_3__22, 
         linha4_3__21, linha4_3__20, linha4_3__19, linha4_3__18, linha4_3__17, 
         linha4_3__16, linha4_3__15, linha4_3__14, linha4_3__13, linha4_3__12, 
         linha4_3__11, linha4_3__10, linha4_3__9, linha4_3__8, linha4_3__7, 
         linha4_3__6, linha4_3__5, linha4_3__4, linha4_3__3, linha4_3__2, 
         linha4_3__1, linha4_3__0, linha4_2__31, linha4_2__30, linha4_2__29, 
         linha4_2__28, linha4_2__27, linha4_2__26, linha4_2__25, linha4_2__24, 
         linha4_2__23, linha4_2__22, linha4_2__21, linha4_2__20, linha4_2__19, 
         linha4_2__18, linha4_2__17, linha4_2__16, linha4_2__15, linha4_2__14, 
         linha4_2__13, linha4_2__12, linha4_2__11, linha4_2__10, linha4_2__9, 
         linha4_2__8, linha4_2__7, linha4_2__6, linha4_2__5, linha4_2__4, 
         linha4_2__3, linha4_2__2, linha4_2__1, linha4_2__0, linha4_1__31, 
         linha4_1__30, linha4_1__29, linha4_1__28, linha4_1__27, linha4_1__26, 
         linha4_1__25, linha4_1__24, linha4_1__23, linha4_1__22, linha4_1__21, 
         linha4_1__20, linha4_1__19, linha4_1__18, linha4_1__17, linha4_1__16, 
         linha4_1__15, linha4_1__14, linha4_1__13, linha4_1__12, linha4_1__11, 
         linha4_1__10, linha4_1__9, linha4_1__8, linha4_1__7, linha4_1__6, 
         linha4_1__5, linha4_1__4, linha4_1__3, linha4_1__2, linha4_1__1, 
         linha4_1__0, linha3_7__31, linha3_7__30, linha3_7__29, linha3_7__28, 
         linha3_7__27, linha3_7__26, linha3_7__25, linha3_7__24, linha3_7__23, 
         linha3_7__22, linha3_7__21, linha3_7__20, linha3_7__19, linha3_7__18, 
         linha3_7__17, linha3_7__16, linha3_7__15, linha3_7__14, linha3_7__13, 
         linha3_7__12, linha3_7__11, linha3_7__10, linha3_7__9, linha3_7__8, 
         linha3_7__7, linha3_7__6, linha3_7__5, linha3_7__4, linha3_7__3, 
         linha3_7__2, linha3_7__1, linha3_7__0, linha3_6__31, linha3_6__30, 
         linha3_6__29, linha3_6__28, linha3_6__27, linha3_6__26, linha3_6__25, 
         linha3_6__24, linha3_6__23, linha3_6__22, linha3_6__21, linha3_6__20, 
         linha3_6__19, linha3_6__18, linha3_6__17, linha3_6__16, linha3_6__15, 
         linha3_6__14, linha3_6__13, linha3_6__12, linha3_6__11, linha3_6__10, 
         linha3_6__9, linha3_6__8, linha3_6__7, linha3_6__6, linha3_6__5, 
         linha3_6__4, linha3_6__3, linha3_6__2, linha3_6__1, linha3_6__0, 
         linha3_5__31, linha3_5__30, linha3_5__29, linha3_5__28, linha3_5__27, 
         linha3_5__26, linha3_5__25, linha3_5__24, linha3_5__23, linha3_5__22, 
         linha3_5__21, linha3_5__20, linha3_5__19, linha3_5__18, linha3_5__17, 
         linha3_5__16, linha3_5__15, linha3_5__14, linha3_5__13, linha3_5__12, 
         linha3_5__11, linha3_5__10, linha3_5__9, linha3_5__8, linha3_5__7, 
         linha3_5__6, linha3_5__5, linha3_5__4, linha3_5__3, linha3_5__2, 
         linha3_5__1, linha3_5__0, linha3_4__31, linha3_4__30, linha3_4__29, 
         linha3_4__28, linha3_4__27, linha3_4__26, linha3_4__25, linha3_4__24, 
         linha3_4__23, linha3_4__22, linha3_4__21, linha3_4__20, linha3_4__19, 
         linha3_4__18, linha3_4__17, linha3_4__16, linha3_4__15, linha3_4__14, 
         linha3_4__13, linha3_4__12, linha3_4__11, linha3_4__10, linha3_4__9, 
         linha3_4__8, linha3_4__7, linha3_4__6, linha3_4__5, linha3_4__4, 
         linha3_4__3, linha3_4__2, linha3_4__1, linha3_4__0, linha3_3__31, 
         linha3_3__30, linha3_3__29, linha3_3__28, linha3_3__27, linha3_3__26, 
         linha3_3__25, linha3_3__24, linha3_3__23, linha3_3__22, linha3_3__21, 
         linha3_3__20, linha3_3__19, linha3_3__18, linha3_3__17, linha3_3__16, 
         linha3_3__15, linha3_3__14, linha3_3__13, linha3_3__12, linha3_3__11, 
         linha3_3__10, linha3_3__9, linha3_3__8, linha3_3__7, linha3_3__6, 
         linha3_3__5, linha3_3__4, linha3_3__3, linha3_3__2, linha3_3__1, 
         linha3_3__0, linha3_2__31, linha3_2__30, linha3_2__29, linha3_2__28, 
         linha3_2__27, linha3_2__26, linha3_2__25, linha3_2__24, linha3_2__23, 
         linha3_2__22, linha3_2__21, linha3_2__20, linha3_2__19, linha3_2__18, 
         linha3_2__17, linha3_2__16, linha3_2__15, linha3_2__14, linha3_2__13, 
         linha3_2__12, linha3_2__11, linha3_2__10, linha3_2__9, linha3_2__8, 
         linha3_2__7, linha3_2__6, linha3_2__5, linha3_2__4, linha3_2__3, 
         linha3_2__2, linha3_2__1, linha3_2__0, linha3_1__31, linha3_1__30, 
         linha3_1__29, linha3_1__28, linha3_1__27, linha3_1__26, linha3_1__25, 
         linha3_1__24, linha3_1__23, linha3_1__22, linha3_1__21, linha3_1__20, 
         linha3_1__19, linha3_1__18, linha3_1__17, linha3_1__16, linha3_1__15, 
         linha3_1__14, linha3_1__13, linha3_1__12, linha3_1__11, linha3_1__10, 
         linha3_1__9, linha3_1__8, linha3_1__7, linha3_1__6, linha3_1__5, 
         linha3_1__4, linha3_1__3, linha3_1__2, linha3_1__1, linha3_1__0, 
         linha2_7__31, linha2_7__30, linha2_7__29, linha2_7__28, linha2_7__27, 
         linha2_7__26, linha2_7__25, linha2_7__24, linha2_7__23, linha2_7__22, 
         linha2_7__21, linha2_7__20, linha2_7__19, linha2_7__18, linha2_7__17, 
         linha2_7__16, linha2_7__15, linha2_7__14, linha2_7__13, linha2_7__12, 
         linha2_7__11, linha2_7__10, linha2_7__9, linha2_7__8, linha2_7__7, 
         linha2_7__6, linha2_7__5, linha2_7__4, linha2_7__3, linha2_7__2, 
         linha2_7__1, linha2_7__0, linha2_6__31, linha2_6__30, linha2_6__29, 
         linha2_6__28, linha2_6__27, linha2_6__26, linha2_6__25, linha2_6__24, 
         linha2_6__23, linha2_6__22, linha2_6__21, linha2_6__20, linha2_6__19, 
         linha2_6__18, linha2_6__17, linha2_6__16, linha2_6__15, linha2_6__14, 
         linha2_6__13, linha2_6__12, linha2_6__11, linha2_6__10, linha2_6__9, 
         linha2_6__8, linha2_6__7, linha2_6__6, linha2_6__5, linha2_6__4, 
         linha2_6__3, linha2_6__2, linha2_6__1, linha2_6__0, linha2_5__31, 
         linha2_5__30, linha2_5__29, linha2_5__28, linha2_5__27, linha2_5__26, 
         linha2_5__25, linha2_5__24, linha2_5__23, linha2_5__22, linha2_5__21, 
         linha2_5__20, linha2_5__19, linha2_5__18, linha2_5__17, linha2_5__16, 
         linha2_5__15, linha2_5__14, linha2_5__13, linha2_5__12, linha2_5__11, 
         linha2_5__10, linha2_5__9, linha2_5__8, linha2_5__7, linha2_5__6, 
         linha2_5__5, linha2_5__4, linha2_5__3, linha2_5__2, linha2_5__1, 
         linha2_5__0, linha2_4__31, linha2_4__30, linha2_4__29, linha2_4__28, 
         linha2_4__27, linha2_4__26, linha2_4__25, linha2_4__24, linha2_4__23, 
         linha2_4__22, linha2_4__21, linha2_4__20, linha2_4__19, linha2_4__18, 
         linha2_4__17, linha2_4__16, linha2_4__15, linha2_4__14, linha2_4__13, 
         linha2_4__12, linha2_4__11, linha2_4__10, linha2_4__9, linha2_4__8, 
         linha2_4__7, linha2_4__6, linha2_4__5, linha2_4__4, linha2_4__3, 
         linha2_4__2, linha2_4__1, linha2_4__0, linha2_3__31, linha2_3__30, 
         linha2_3__29, linha2_3__28, linha2_3__27, linha2_3__26, linha2_3__25, 
         linha2_3__24, linha2_3__23, linha2_3__22, linha2_3__21, linha2_3__20, 
         linha2_3__19, linha2_3__18, linha2_3__17, linha2_3__16, linha2_3__15, 
         linha2_3__14, linha2_3__13, linha2_3__12, linha2_3__11, linha2_3__10, 
         linha2_3__9, linha2_3__8, linha2_3__7, linha2_3__6, linha2_3__5, 
         linha2_3__4, linha2_3__3, linha2_3__2, linha2_3__1, linha2_3__0, 
         linha2_2__31, linha2_2__30, linha2_2__29, linha2_2__28, linha2_2__27, 
         linha2_2__26, linha2_2__25, linha2_2__24, linha2_2__23, linha2_2__22, 
         linha2_2__21, linha2_2__20, linha2_2__19, linha2_2__18, linha2_2__17, 
         linha2_2__16, linha2_2__15, linha2_2__14, linha2_2__13, linha2_2__12, 
         linha2_2__11, linha2_2__10, linha2_2__9, linha2_2__8, linha2_2__7, 
         linha2_2__6, linha2_2__5, linha2_2__4, linha2_2__3, linha2_2__2, 
         linha2_2__1, linha2_2__0, linha2_1__31, linha2_1__30, linha2_1__29, 
         linha2_1__28, linha2_1__27, linha2_1__26, linha2_1__25, linha2_1__24, 
         linha2_1__23, linha2_1__22, linha2_1__21, linha2_1__20, linha2_1__19, 
         linha2_1__18, linha2_1__17, linha2_1__16, linha2_1__15, linha2_1__14, 
         linha2_1__13, linha2_1__12, linha2_1__11, linha2_1__10, linha2_1__9, 
         linha2_1__8, linha2_1__7, linha2_1__6, linha2_1__5, linha2_1__4, 
         linha2_1__3, linha2_1__2, linha2_1__1, linha2_1__0, linha8_3__31, 
         linha8_3__30, linha8_3__29, linha8_3__28, linha8_3__27, linha8_3__26, 
         linha8_3__25, linha8_3__24, linha8_3__23, linha8_3__22, linha8_3__21, 
         linha8_3__20, linha8_3__19, linha8_3__18, linha8_3__17, linha8_3__16, 
         linha8_3__15, linha8_3__14, linha8_3__13, linha8_3__12, linha8_3__11, 
         linha8_3__10, linha8_3__9, linha8_3__8, linha8_3__7, linha8_3__6, 
         linha8_3__5, linha8_3__4, linha8_3__3, linha8_3__2, linha8_3__1, 
         linha8_3__0, linha8_2__31, linha8_2__30, linha8_2__29, linha8_2__28, 
         linha8_2__27, linha8_2__26, linha8_2__25, linha8_2__24, linha8_2__23, 
         linha8_2__22, linha8_2__21, linha8_2__20, linha8_2__19, linha8_2__18, 
         linha8_2__17, linha8_2__16, linha8_2__15, linha8_2__14, linha8_2__13, 
         linha8_2__12, linha8_2__11, linha8_2__10, linha8_2__9, linha8_2__8, 
         linha8_2__7, linha8_2__6, linha8_2__5, linha8_2__4, linha8_2__3, 
         linha8_2__2, linha8_2__1, linha8_2__0, linha8_1__31, linha8_1__30, 
         linha8_1__29, linha8_1__28, linha8_1__27, linha8_1__26, linha8_1__25, 
         linha8_1__24, linha8_1__23, linha8_1__22, linha8_1__21, linha8_1__20, 
         linha8_1__19, linha8_1__18, linha8_1__17, linha8_1__16, linha8_1__15, 
         linha8_1__14, linha8_1__13, linha8_1__12, linha8_1__11, linha8_1__10, 
         linha8_1__9, linha8_1__8, linha8_1__7, linha8_1__6, linha8_1__5, 
         linha8_1__4, linha8_1__3, linha8_1__2, linha8_1__1, linha8_1__0, 
         linha1_3__31, linha1_3__30, linha1_3__29, linha1_3__28, linha1_3__27, 
         linha1_3__26, linha1_3__25, linha1_3__24, linha1_3__23, linha1_3__22, 
         linha1_3__21, linha1_3__20, linha1_3__19, linha1_3__18, linha1_3__17, 
         linha1_3__16, linha1_3__15, linha1_3__14, linha1_3__13, linha1_3__12, 
         linha1_3__11, linha1_3__10, linha1_3__9, linha1_3__8, linha1_3__7, 
         linha1_3__6, linha1_3__5, linha1_3__4, linha1_3__3, linha1_3__2, 
         linha1_3__1, linha1_3__0, linha1_2__31, linha1_2__30, linha1_2__29, 
         linha1_2__28, linha1_2__27, linha1_2__26, linha1_2__25, linha1_2__24, 
         linha1_2__23, linha1_2__22, linha1_2__21, linha1_2__20, linha1_2__19, 
         linha1_2__18, linha1_2__17, linha1_2__16, linha1_2__15, linha1_2__14, 
         linha1_2__13, linha1_2__12, linha1_2__11, linha1_2__10, linha1_2__9, 
         linha1_2__8, linha1_2__7, linha1_2__6, linha1_2__5, linha1_2__4, 
         linha1_2__3, linha1_2__2, linha1_2__1, linha1_2__0, linha1_1__31, 
         linha1_1__30, linha1_1__29, linha1_1__28, linha1_1__27, linha1_1__26, 
         linha1_1__25, linha1_1__24, linha1_1__23, linha1_1__22, linha1_1__21, 
         linha1_1__20, linha1_1__19, linha1_1__18, linha1_1__17, linha1_1__16, 
         linha1_1__15, linha1_1__14, linha1_1__13, linha1_1__12, linha1_1__11, 
         linha1_1__10, linha1_1__9, linha1_1__8, linha1_1__7, linha1_1__6, 
         linha1_1__5, linha1_1__4, linha1_1__3, linha1_1__2, linha1_1__1, 
         linha1_1__0, row_0_rowp_bni1_l, row_0_rowp_bni2_l, row_0_rowp_bni3_l, 
         row_0_rowp_bni4_l, row_1_rowi_bni1_l, row_1_rowi_bni2_l, 
         row_1_rowi_bni3_l, row_2_rowp_bni1_l, row_2_rowp_bni2_l, 
         row_2_rowp_bni3_l, row_2_rowp_bni4_l, row_3_rowi_bni1_l, 
         row_3_rowi_bni2_l, row_3_rowi_bni3_l, row_4_rowp_bni1_l, 
         row_4_rowp_bni2_l, row_4_rowp_bni3_l, row_4_rowp_bni4_l, 
         row_5_rowi_bni1_l, row_5_rowi_bni2_l, row_5_rowi_bni3_l, 
         row_6_rowp_bni1_l, row_6_rowp_bni2_l, row_6_rowp_bni3_l, 
         row_6_rowp_bni4_l, row_7_rowi_bni1_l, row_7_rowi_bni2_l, 
         row_7_rowi_bni3_l, nx4095;
    wire [27:0] \$dummy ;




    juntarComparadores_32 row_0_rowp_bni1_Comp (.g (\$dummy [0]), .l (
                          row_0_rowp_bni1_l), .a ({x1[31],x1[30],x1[29],x1[28],
                          x1[27],x1[26],x1[25],x1[24],x1[23],x1[22],x1[21],
                          x1[20],x1[19],x1[18],x1[17],x1[16],x1[15],x1[14],
                          x1[13],x1[12],x1[11],x1[10],x1[9],x1[8],x1[7],x1[6],
                          x1[5],x1[4],x1[3],x1[2],x1[1],x1[0]}), .b ({x2[31],
                          x2[30],x2[29],x2[28],x2[27],x2[26],x2[25],x2[24],
                          x2[23],x2[22],x2[21],x2[20],x2[19],x2[18],x2[17],
                          x2[16],x2[15],x2[14],x2[13],x2[12],x2[11],x2[10],x2[9]
                          ,x2[8],x2[7],x2[6],x2[5],x2[4],x2[3],x2[2],x2[1],x2[0]
                          })) ;
    Mux2x1_32 row_0_rowp_bni1_muxMax (.r ({linha1_1__31,linha1_1__30,
              linha1_1__29,linha1_1__28,linha1_1__27,linha1_1__26,linha1_1__25,
              linha1_1__24,linha1_1__23,linha1_1__22,linha1_1__21,linha1_1__20,
              linha1_1__19,linha1_1__18,linha1_1__17,linha1_1__16,linha1_1__15,
              linha1_1__14,linha1_1__13,linha1_1__12,linha1_1__11,linha1_1__10,
              linha1_1__9,linha1_1__8,linha1_1__7,linha1_1__6,linha1_1__5,
              linha1_1__4,linha1_1__3,linha1_1__2,linha1_1__1,linha1_1__0}), .a1 (
              {x2[31],x2[30],x2[29],x2[28],x2[27],x2[26],x2[25],x2[24],x2[23],
              x2[22],x2[21],x2[20],x2[19],x2[18],x2[17],x2[16],x2[15],x2[14],
              x2[13],x2[12],x2[11],x2[10],x2[9],x2[8],x2[7],x2[6],x2[5],x2[4],
              x2[3],x2[2],x2[1],x2[0]}), .a0 ({x1[31],x1[30],x1[29],x1[28],
              x1[27],x1[26],x1[25],x1[24],x1[23],x1[22],x1[21],x1[20],x1[19],
              x1[18],x1[17],x1[16],x1[15],x1[14],x1[13],x1[12],x1[11],x1[10],
              x1[9],x1[8],x1[7],x1[6],x1[5],x1[4],x1[3],x1[2],x1[1],x1[0]}), .s (
              nx4095)) ;
    Mux2x1_32 row_0_rowp_bni1_muxMin (.r ({linha2_1__31,linha2_1__30,
              linha2_1__29,linha2_1__28,linha2_1__27,linha2_1__26,linha2_1__25,
              linha2_1__24,linha2_1__23,linha2_1__22,linha2_1__21,linha2_1__20,
              linha2_1__19,linha2_1__18,linha2_1__17,linha2_1__16,linha2_1__15,
              linha2_1__14,linha2_1__13,linha2_1__12,linha2_1__11,linha2_1__10,
              linha2_1__9,linha2_1__8,linha2_1__7,linha2_1__6,linha2_1__5,
              linha2_1__4,linha2_1__3,linha2_1__2,linha2_1__1,linha2_1__0}), .a1 (
              {x1[31],x1[30],x1[29],x1[28],x1[27],x1[26],x1[25],x1[24],x1[23],
              x1[22],x1[21],x1[20],x1[19],x1[18],x1[17],x1[16],x1[15],x1[14],
              x1[13],x1[12],x1[11],x1[10],x1[9],x1[8],x1[7],x1[6],x1[5],x1[4],
              x1[3],x1[2],x1[1],x1[0]}), .a0 ({x2[31],x2[30],x2[29],x2[28],
              x2[27],x2[26],x2[25],x2[24],x2[23],x2[22],x2[21],x2[20],x2[19],
              x2[18],x2[17],x2[16],x2[15],x2[14],x2[13],x2[12],x2[11],x2[10],
              x2[9],x2[8],x2[7],x2[6],x2[5],x2[4],x2[3],x2[2],x2[1],x2[0]}), .s (
              nx4095)) ;
    juntarComparadores_32 row_0_rowp_bni2_Comp (.g (\$dummy [1]), .l (
                          row_0_rowp_bni2_l), .a ({x3[31],x3[30],x3[29],x3[28],
                          x3[27],x3[26],x3[25],x3[24],x3[23],x3[22],x3[21],
                          x3[20],x3[19],x3[18],x3[17],x3[16],x3[15],x3[14],
                          x3[13],x3[12],x3[11],x3[10],x3[9],x3[8],x3[7],x3[6],
                          x3[5],x3[4],x3[3],x3[2],x3[1],x3[0]}), .b ({x4[31],
                          x4[30],x4[29],x4[28],x4[27],x4[26],x4[25],x4[24],
                          x4[23],x4[22],x4[21],x4[20],x4[19],x4[18],x4[17],
                          x4[16],x4[15],x4[14],x4[13],x4[12],x4[11],x4[10],x4[9]
                          ,x4[8],x4[7],x4[6],x4[5],x4[4],x4[3],x4[2],x4[1],x4[0]
                          })) ;
    Mux2x1_32 row_0_rowp_bni2_muxMax (.r ({linha3_1__31,linha3_1__30,
              linha3_1__29,linha3_1__28,linha3_1__27,linha3_1__26,linha3_1__25,
              linha3_1__24,linha3_1__23,linha3_1__22,linha3_1__21,linha3_1__20,
              linha3_1__19,linha3_1__18,linha3_1__17,linha3_1__16,linha3_1__15,
              linha3_1__14,linha3_1__13,linha3_1__12,linha3_1__11,linha3_1__10,
              linha3_1__9,linha3_1__8,linha3_1__7,linha3_1__6,linha3_1__5,
              linha3_1__4,linha3_1__3,linha3_1__2,linha3_1__1,linha3_1__0}), .a1 (
              {x4[31],x4[30],x4[29],x4[28],x4[27],x4[26],x4[25],x4[24],x4[23],
              x4[22],x4[21],x4[20],x4[19],x4[18],x4[17],x4[16],x4[15],x4[14],
              x4[13],x4[12],x4[11],x4[10],x4[9],x4[8],x4[7],x4[6],x4[5],x4[4],
              x4[3],x4[2],x4[1],x4[0]}), .a0 ({x3[31],x3[30],x3[29],x3[28],
              x3[27],x3[26],x3[25],x3[24],x3[23],x3[22],x3[21],x3[20],x3[19],
              x3[18],x3[17],x3[16],x3[15],x3[14],x3[13],x3[12],x3[11],x3[10],
              x3[9],x3[8],x3[7],x3[6],x3[5],x3[4],x3[3],x3[2],x3[1],x3[0]}), .s (
              row_0_rowp_bni2_l)) ;
    Mux2x1_32 row_0_rowp_bni2_muxMin (.r ({linha4_1__31,linha4_1__30,
              linha4_1__29,linha4_1__28,linha4_1__27,linha4_1__26,linha4_1__25,
              linha4_1__24,linha4_1__23,linha4_1__22,linha4_1__21,linha4_1__20,
              linha4_1__19,linha4_1__18,linha4_1__17,linha4_1__16,linha4_1__15,
              linha4_1__14,linha4_1__13,linha4_1__12,linha4_1__11,linha4_1__10,
              linha4_1__9,linha4_1__8,linha4_1__7,linha4_1__6,linha4_1__5,
              linha4_1__4,linha4_1__3,linha4_1__2,linha4_1__1,linha4_1__0}), .a1 (
              {x3[31],x3[30],x3[29],x3[28],x3[27],x3[26],x3[25],x3[24],x3[23],
              x3[22],x3[21],x3[20],x3[19],x3[18],x3[17],x3[16],x3[15],x3[14],
              x3[13],x3[12],x3[11],x3[10],x3[9],x3[8],x3[7],x3[6],x3[5],x3[4],
              x3[3],x3[2],x3[1],x3[0]}), .a0 ({x4[31],x4[30],x4[29],x4[28],
              x4[27],x4[26],x4[25],x4[24],x4[23],x4[22],x4[21],x4[20],x4[19],
              x4[18],x4[17],x4[16],x4[15],x4[14],x4[13],x4[12],x4[11],x4[10],
              x4[9],x4[8],x4[7],x4[6],x4[5],x4[4],x4[3],x4[2],x4[1],x4[0]}), .s (
              row_0_rowp_bni2_l)) ;
    juntarComparadores_32 row_0_rowp_bni3_Comp (.g (\$dummy [2]), .l (
                          row_0_rowp_bni3_l), .a ({x5[31],x5[30],x5[29],x5[28],
                          x5[27],x5[26],x5[25],x5[24],x5[23],x5[22],x5[21],
                          x5[20],x5[19],x5[18],x5[17],x5[16],x5[15],x5[14],
                          x5[13],x5[12],x5[11],x5[10],x5[9],x5[8],x5[7],x5[6],
                          x5[5],x5[4],x5[3],x5[2],x5[1],x5[0]}), .b ({x6[31],
                          x6[30],x6[29],x6[28],x6[27],x6[26],x6[25],x6[24],
                          x6[23],x6[22],x6[21],x6[20],x6[19],x6[18],x6[17],
                          x6[16],x6[15],x6[14],x6[13],x6[12],x6[11],x6[10],x6[9]
                          ,x6[8],x6[7],x6[6],x6[5],x6[4],x6[3],x6[2],x6[1],x6[0]
                          })) ;
    Mux2x1_32 row_0_rowp_bni3_muxMax (.r ({linha5_1__31,linha5_1__30,
              linha5_1__29,linha5_1__28,linha5_1__27,linha5_1__26,linha5_1__25,
              linha5_1__24,linha5_1__23,linha5_1__22,linha5_1__21,linha5_1__20,
              linha5_1__19,linha5_1__18,linha5_1__17,linha5_1__16,linha5_1__15,
              linha5_1__14,linha5_1__13,linha5_1__12,linha5_1__11,linha5_1__10,
              linha5_1__9,linha5_1__8,linha5_1__7,linha5_1__6,linha5_1__5,
              linha5_1__4,linha5_1__3,linha5_1__2,linha5_1__1,linha5_1__0}), .a1 (
              {x6[31],x6[30],x6[29],x6[28],x6[27],x6[26],x6[25],x6[24],x6[23],
              x6[22],x6[21],x6[20],x6[19],x6[18],x6[17],x6[16],x6[15],x6[14],
              x6[13],x6[12],x6[11],x6[10],x6[9],x6[8],x6[7],x6[6],x6[5],x6[4],
              x6[3],x6[2],x6[1],x6[0]}), .a0 ({x5[31],x5[30],x5[29],x5[28],
              x5[27],x5[26],x5[25],x5[24],x5[23],x5[22],x5[21],x5[20],x5[19],
              x5[18],x5[17],x5[16],x5[15],x5[14],x5[13],x5[12],x5[11],x5[10],
              x5[9],x5[8],x5[7],x5[6],x5[5],x5[4],x5[3],x5[2],x5[1],x5[0]}), .s (
              row_0_rowp_bni3_l)) ;
    Mux2x1_32 row_0_rowp_bni3_muxMin (.r ({linha6_1__31,linha6_1__30,
              linha6_1__29,linha6_1__28,linha6_1__27,linha6_1__26,linha6_1__25,
              linha6_1__24,linha6_1__23,linha6_1__22,linha6_1__21,linha6_1__20,
              linha6_1__19,linha6_1__18,linha6_1__17,linha6_1__16,linha6_1__15,
              linha6_1__14,linha6_1__13,linha6_1__12,linha6_1__11,linha6_1__10,
              linha6_1__9,linha6_1__8,linha6_1__7,linha6_1__6,linha6_1__5,
              linha6_1__4,linha6_1__3,linha6_1__2,linha6_1__1,linha6_1__0}), .a1 (
              {x5[31],x5[30],x5[29],x5[28],x5[27],x5[26],x5[25],x5[24],x5[23],
              x5[22],x5[21],x5[20],x5[19],x5[18],x5[17],x5[16],x5[15],x5[14],
              x5[13],x5[12],x5[11],x5[10],x5[9],x5[8],x5[7],x5[6],x5[5],x5[4],
              x5[3],x5[2],x5[1],x5[0]}), .a0 ({x6[31],x6[30],x6[29],x6[28],
              x6[27],x6[26],x6[25],x6[24],x6[23],x6[22],x6[21],x6[20],x6[19],
              x6[18],x6[17],x6[16],x6[15],x6[14],x6[13],x6[12],x6[11],x6[10],
              x6[9],x6[8],x6[7],x6[6],x6[5],x6[4],x6[3],x6[2],x6[1],x6[0]}), .s (
              row_0_rowp_bni3_l)) ;
    juntarComparadores_32 row_0_rowp_bni4_Comp (.g (\$dummy [3]), .l (
                          row_0_rowp_bni4_l), .a ({x7[31],x7[30],x7[29],x7[28],
                          x7[27],x7[26],x7[25],x7[24],x7[23],x7[22],x7[21],
                          x7[20],x7[19],x7[18],x7[17],x7[16],x7[15],x7[14],
                          x7[13],x7[12],x7[11],x7[10],x7[9],x7[8],x7[7],x7[6],
                          x7[5],x7[4],x7[3],x7[2],x7[1],x7[0]}), .b ({x8[31],
                          x8[30],x8[29],x8[28],x8[27],x8[26],x8[25],x8[24],
                          x8[23],x8[22],x8[21],x8[20],x8[19],x8[18],x8[17],
                          x8[16],x8[15],x8[14],x8[13],x8[12],x8[11],x8[10],x8[9]
                          ,x8[8],x8[7],x8[6],x8[5],x8[4],x8[3],x8[2],x8[1],x8[0]
                          })) ;
    Mux2x1_32 row_0_rowp_bni4_muxMax (.r ({linha7_1__31,linha7_1__30,
              linha7_1__29,linha7_1__28,linha7_1__27,linha7_1__26,linha7_1__25,
              linha7_1__24,linha7_1__23,linha7_1__22,linha7_1__21,linha7_1__20,
              linha7_1__19,linha7_1__18,linha7_1__17,linha7_1__16,linha7_1__15,
              linha7_1__14,linha7_1__13,linha7_1__12,linha7_1__11,linha7_1__10,
              linha7_1__9,linha7_1__8,linha7_1__7,linha7_1__6,linha7_1__5,
              linha7_1__4,linha7_1__3,linha7_1__2,linha7_1__1,linha7_1__0}), .a1 (
              {x8[31],x8[30],x8[29],x8[28],x8[27],x8[26],x8[25],x8[24],x8[23],
              x8[22],x8[21],x8[20],x8[19],x8[18],x8[17],x8[16],x8[15],x8[14],
              x8[13],x8[12],x8[11],x8[10],x8[9],x8[8],x8[7],x8[6],x8[5],x8[4],
              x8[3],x8[2],x8[1],x8[0]}), .a0 ({x7[31],x7[30],x7[29],x7[28],
              x7[27],x7[26],x7[25],x7[24],x7[23],x7[22],x7[21],x7[20],x7[19],
              x7[18],x7[17],x7[16],x7[15],x7[14],x7[13],x7[12],x7[11],x7[10],
              x7[9],x7[8],x7[7],x7[6],x7[5],x7[4],x7[3],x7[2],x7[1],x7[0]}), .s (
              row_0_rowp_bni4_l)) ;
    Mux2x1_32 row_0_rowp_bni4_muxMin (.r ({linha8_1__31,linha8_1__30,
              linha8_1__29,linha8_1__28,linha8_1__27,linha8_1__26,linha8_1__25,
              linha8_1__24,linha8_1__23,linha8_1__22,linha8_1__21,linha8_1__20,
              linha8_1__19,linha8_1__18,linha8_1__17,linha8_1__16,linha8_1__15,
              linha8_1__14,linha8_1__13,linha8_1__12,linha8_1__11,linha8_1__10,
              linha8_1__9,linha8_1__8,linha8_1__7,linha8_1__6,linha8_1__5,
              linha8_1__4,linha8_1__3,linha8_1__2,linha8_1__1,linha8_1__0}), .a1 (
              {x7[31],x7[30],x7[29],x7[28],x7[27],x7[26],x7[25],x7[24],x7[23],
              x7[22],x7[21],x7[20],x7[19],x7[18],x7[17],x7[16],x7[15],x7[14],
              x7[13],x7[12],x7[11],x7[10],x7[9],x7[8],x7[7],x7[6],x7[5],x7[4],
              x7[3],x7[2],x7[1],x7[0]}), .a0 ({x8[31],x8[30],x8[29],x8[28],
              x8[27],x8[26],x8[25],x8[24],x8[23],x8[22],x8[21],x8[20],x8[19],
              x8[18],x8[17],x8[16],x8[15],x8[14],x8[13],x8[12],x8[11],x8[10],
              x8[9],x8[8],x8[7],x8[6],x8[5],x8[4],x8[3],x8[2],x8[1],x8[0]}), .s (
              row_0_rowp_bni4_l)) ;
    juntarComparadores_32 row_1_rowi_bni1_Comp (.g (\$dummy [4]), .l (
                          row_1_rowi_bni1_l), .a ({linha2_1__31,linha2_1__30,
                          linha2_1__29,linha2_1__28,linha2_1__27,linha2_1__26,
                          linha2_1__25,linha2_1__24,linha2_1__23,linha2_1__22,
                          linha2_1__21,linha2_1__20,linha2_1__19,linha2_1__18,
                          linha2_1__17,linha2_1__16,linha2_1__15,linha2_1__14,
                          linha2_1__13,linha2_1__12,linha2_1__11,linha2_1__10,
                          linha2_1__9,linha2_1__8,linha2_1__7,linha2_1__6,
                          linha2_1__5,linha2_1__4,linha2_1__3,linha2_1__2,
                          linha2_1__1,linha2_1__0}), .b ({linha3_1__31,
                          linha3_1__30,linha3_1__29,linha3_1__28,linha3_1__27,
                          linha3_1__26,linha3_1__25,linha3_1__24,linha3_1__23,
                          linha3_1__22,linha3_1__21,linha3_1__20,linha3_1__19,
                          linha3_1__18,linha3_1__17,linha3_1__16,linha3_1__15,
                          linha3_1__14,linha3_1__13,linha3_1__12,linha3_1__11,
                          linha3_1__10,linha3_1__9,linha3_1__8,linha3_1__7,
                          linha3_1__6,linha3_1__5,linha3_1__4,linha3_1__3,
                          linha3_1__2,linha3_1__1,linha3_1__0})) ;
    Mux2x1_32 row_1_rowi_bni1_muxMax (.r ({linha2_2__31,linha2_2__30,
              linha2_2__29,linha2_2__28,linha2_2__27,linha2_2__26,linha2_2__25,
              linha2_2__24,linha2_2__23,linha2_2__22,linha2_2__21,linha2_2__20,
              linha2_2__19,linha2_2__18,linha2_2__17,linha2_2__16,linha2_2__15,
              linha2_2__14,linha2_2__13,linha2_2__12,linha2_2__11,linha2_2__10,
              linha2_2__9,linha2_2__8,linha2_2__7,linha2_2__6,linha2_2__5,
              linha2_2__4,linha2_2__3,linha2_2__2,linha2_2__1,linha2_2__0}), .a1 (
              {linha3_1__31,linha3_1__30,linha3_1__29,linha3_1__28,linha3_1__27,
              linha3_1__26,linha3_1__25,linha3_1__24,linha3_1__23,linha3_1__22,
              linha3_1__21,linha3_1__20,linha3_1__19,linha3_1__18,linha3_1__17,
              linha3_1__16,linha3_1__15,linha3_1__14,linha3_1__13,linha3_1__12,
              linha3_1__11,linha3_1__10,linha3_1__9,linha3_1__8,linha3_1__7,
              linha3_1__6,linha3_1__5,linha3_1__4,linha3_1__3,linha3_1__2,
              linha3_1__1,linha3_1__0}), .a0 ({linha2_1__31,linha2_1__30,
              linha2_1__29,linha2_1__28,linha2_1__27,linha2_1__26,linha2_1__25,
              linha2_1__24,linha2_1__23,linha2_1__22,linha2_1__21,linha2_1__20,
              linha2_1__19,linha2_1__18,linha2_1__17,linha2_1__16,linha2_1__15,
              linha2_1__14,linha2_1__13,linha2_1__12,linha2_1__11,linha2_1__10,
              linha2_1__9,linha2_1__8,linha2_1__7,linha2_1__6,linha2_1__5,
              linha2_1__4,linha2_1__3,linha2_1__2,linha2_1__1,linha2_1__0}), .s (
              row_1_rowi_bni1_l)) ;
    Mux2x1_32 row_1_rowi_bni1_muxMin (.r ({linha3_2__31,linha3_2__30,
              linha3_2__29,linha3_2__28,linha3_2__27,linha3_2__26,linha3_2__25,
              linha3_2__24,linha3_2__23,linha3_2__22,linha3_2__21,linha3_2__20,
              linha3_2__19,linha3_2__18,linha3_2__17,linha3_2__16,linha3_2__15,
              linha3_2__14,linha3_2__13,linha3_2__12,linha3_2__11,linha3_2__10,
              linha3_2__9,linha3_2__8,linha3_2__7,linha3_2__6,linha3_2__5,
              linha3_2__4,linha3_2__3,linha3_2__2,linha3_2__1,linha3_2__0}), .a1 (
              {linha2_1__31,linha2_1__30,linha2_1__29,linha2_1__28,linha2_1__27,
              linha2_1__26,linha2_1__25,linha2_1__24,linha2_1__23,linha2_1__22,
              linha2_1__21,linha2_1__20,linha2_1__19,linha2_1__18,linha2_1__17,
              linha2_1__16,linha2_1__15,linha2_1__14,linha2_1__13,linha2_1__12,
              linha2_1__11,linha2_1__10,linha2_1__9,linha2_1__8,linha2_1__7,
              linha2_1__6,linha2_1__5,linha2_1__4,linha2_1__3,linha2_1__2,
              linha2_1__1,linha2_1__0}), .a0 ({linha3_1__31,linha3_1__30,
              linha3_1__29,linha3_1__28,linha3_1__27,linha3_1__26,linha3_1__25,
              linha3_1__24,linha3_1__23,linha3_1__22,linha3_1__21,linha3_1__20,
              linha3_1__19,linha3_1__18,linha3_1__17,linha3_1__16,linha3_1__15,
              linha3_1__14,linha3_1__13,linha3_1__12,linha3_1__11,linha3_1__10,
              linha3_1__9,linha3_1__8,linha3_1__7,linha3_1__6,linha3_1__5,
              linha3_1__4,linha3_1__3,linha3_1__2,linha3_1__1,linha3_1__0}), .s (
              row_1_rowi_bni1_l)) ;
    juntarComparadores_32 row_1_rowi_bni2_Comp (.g (\$dummy [5]), .l (
                          row_1_rowi_bni2_l), .a ({linha4_1__31,linha4_1__30,
                          linha4_1__29,linha4_1__28,linha4_1__27,linha4_1__26,
                          linha4_1__25,linha4_1__24,linha4_1__23,linha4_1__22,
                          linha4_1__21,linha4_1__20,linha4_1__19,linha4_1__18,
                          linha4_1__17,linha4_1__16,linha4_1__15,linha4_1__14,
                          linha4_1__13,linha4_1__12,linha4_1__11,linha4_1__10,
                          linha4_1__9,linha4_1__8,linha4_1__7,linha4_1__6,
                          linha4_1__5,linha4_1__4,linha4_1__3,linha4_1__2,
                          linha4_1__1,linha4_1__0}), .b ({linha5_1__31,
                          linha5_1__30,linha5_1__29,linha5_1__28,linha5_1__27,
                          linha5_1__26,linha5_1__25,linha5_1__24,linha5_1__23,
                          linha5_1__22,linha5_1__21,linha5_1__20,linha5_1__19,
                          linha5_1__18,linha5_1__17,linha5_1__16,linha5_1__15,
                          linha5_1__14,linha5_1__13,linha5_1__12,linha5_1__11,
                          linha5_1__10,linha5_1__9,linha5_1__8,linha5_1__7,
                          linha5_1__6,linha5_1__5,linha5_1__4,linha5_1__3,
                          linha5_1__2,linha5_1__1,linha5_1__0})) ;
    Mux2x1_32 row_1_rowi_bni2_muxMax (.r ({linha4_2__31,linha4_2__30,
              linha4_2__29,linha4_2__28,linha4_2__27,linha4_2__26,linha4_2__25,
              linha4_2__24,linha4_2__23,linha4_2__22,linha4_2__21,linha4_2__20,
              linha4_2__19,linha4_2__18,linha4_2__17,linha4_2__16,linha4_2__15,
              linha4_2__14,linha4_2__13,linha4_2__12,linha4_2__11,linha4_2__10,
              linha4_2__9,linha4_2__8,linha4_2__7,linha4_2__6,linha4_2__5,
              linha4_2__4,linha4_2__3,linha4_2__2,linha4_2__1,linha4_2__0}), .a1 (
              {linha5_1__31,linha5_1__30,linha5_1__29,linha5_1__28,linha5_1__27,
              linha5_1__26,linha5_1__25,linha5_1__24,linha5_1__23,linha5_1__22,
              linha5_1__21,linha5_1__20,linha5_1__19,linha5_1__18,linha5_1__17,
              linha5_1__16,linha5_1__15,linha5_1__14,linha5_1__13,linha5_1__12,
              linha5_1__11,linha5_1__10,linha5_1__9,linha5_1__8,linha5_1__7,
              linha5_1__6,linha5_1__5,linha5_1__4,linha5_1__3,linha5_1__2,
              linha5_1__1,linha5_1__0}), .a0 ({linha4_1__31,linha4_1__30,
              linha4_1__29,linha4_1__28,linha4_1__27,linha4_1__26,linha4_1__25,
              linha4_1__24,linha4_1__23,linha4_1__22,linha4_1__21,linha4_1__20,
              linha4_1__19,linha4_1__18,linha4_1__17,linha4_1__16,linha4_1__15,
              linha4_1__14,linha4_1__13,linha4_1__12,linha4_1__11,linha4_1__10,
              linha4_1__9,linha4_1__8,linha4_1__7,linha4_1__6,linha4_1__5,
              linha4_1__4,linha4_1__3,linha4_1__2,linha4_1__1,linha4_1__0}), .s (
              row_1_rowi_bni2_l)) ;
    Mux2x1_32 row_1_rowi_bni2_muxMin (.r ({linha5_2__31,linha5_2__30,
              linha5_2__29,linha5_2__28,linha5_2__27,linha5_2__26,linha5_2__25,
              linha5_2__24,linha5_2__23,linha5_2__22,linha5_2__21,linha5_2__20,
              linha5_2__19,linha5_2__18,linha5_2__17,linha5_2__16,linha5_2__15,
              linha5_2__14,linha5_2__13,linha5_2__12,linha5_2__11,linha5_2__10,
              linha5_2__9,linha5_2__8,linha5_2__7,linha5_2__6,linha5_2__5,
              linha5_2__4,linha5_2__3,linha5_2__2,linha5_2__1,linha5_2__0}), .a1 (
              {linha4_1__31,linha4_1__30,linha4_1__29,linha4_1__28,linha4_1__27,
              linha4_1__26,linha4_1__25,linha4_1__24,linha4_1__23,linha4_1__22,
              linha4_1__21,linha4_1__20,linha4_1__19,linha4_1__18,linha4_1__17,
              linha4_1__16,linha4_1__15,linha4_1__14,linha4_1__13,linha4_1__12,
              linha4_1__11,linha4_1__10,linha4_1__9,linha4_1__8,linha4_1__7,
              linha4_1__6,linha4_1__5,linha4_1__4,linha4_1__3,linha4_1__2,
              linha4_1__1,linha4_1__0}), .a0 ({linha5_1__31,linha5_1__30,
              linha5_1__29,linha5_1__28,linha5_1__27,linha5_1__26,linha5_1__25,
              linha5_1__24,linha5_1__23,linha5_1__22,linha5_1__21,linha5_1__20,
              linha5_1__19,linha5_1__18,linha5_1__17,linha5_1__16,linha5_1__15,
              linha5_1__14,linha5_1__13,linha5_1__12,linha5_1__11,linha5_1__10,
              linha5_1__9,linha5_1__8,linha5_1__7,linha5_1__6,linha5_1__5,
              linha5_1__4,linha5_1__3,linha5_1__2,linha5_1__1,linha5_1__0}), .s (
              row_1_rowi_bni2_l)) ;
    juntarComparadores_32 row_1_rowi_bni3_Comp (.g (\$dummy [6]), .l (
                          row_1_rowi_bni3_l), .a ({linha6_1__31,linha6_1__30,
                          linha6_1__29,linha6_1__28,linha6_1__27,linha6_1__26,
                          linha6_1__25,linha6_1__24,linha6_1__23,linha6_1__22,
                          linha6_1__21,linha6_1__20,linha6_1__19,linha6_1__18,
                          linha6_1__17,linha6_1__16,linha6_1__15,linha6_1__14,
                          linha6_1__13,linha6_1__12,linha6_1__11,linha6_1__10,
                          linha6_1__9,linha6_1__8,linha6_1__7,linha6_1__6,
                          linha6_1__5,linha6_1__4,linha6_1__3,linha6_1__2,
                          linha6_1__1,linha6_1__0}), .b ({linha7_1__31,
                          linha7_1__30,linha7_1__29,linha7_1__28,linha7_1__27,
                          linha7_1__26,linha7_1__25,linha7_1__24,linha7_1__23,
                          linha7_1__22,linha7_1__21,linha7_1__20,linha7_1__19,
                          linha7_1__18,linha7_1__17,linha7_1__16,linha7_1__15,
                          linha7_1__14,linha7_1__13,linha7_1__12,linha7_1__11,
                          linha7_1__10,linha7_1__9,linha7_1__8,linha7_1__7,
                          linha7_1__6,linha7_1__5,linha7_1__4,linha7_1__3,
                          linha7_1__2,linha7_1__1,linha7_1__0})) ;
    Mux2x1_32 row_1_rowi_bni3_muxMax (.r ({linha6_2__31,linha6_2__30,
              linha6_2__29,linha6_2__28,linha6_2__27,linha6_2__26,linha6_2__25,
              linha6_2__24,linha6_2__23,linha6_2__22,linha6_2__21,linha6_2__20,
              linha6_2__19,linha6_2__18,linha6_2__17,linha6_2__16,linha6_2__15,
              linha6_2__14,linha6_2__13,linha6_2__12,linha6_2__11,linha6_2__10,
              linha6_2__9,linha6_2__8,linha6_2__7,linha6_2__6,linha6_2__5,
              linha6_2__4,linha6_2__3,linha6_2__2,linha6_2__1,linha6_2__0}), .a1 (
              {linha7_1__31,linha7_1__30,linha7_1__29,linha7_1__28,linha7_1__27,
              linha7_1__26,linha7_1__25,linha7_1__24,linha7_1__23,linha7_1__22,
              linha7_1__21,linha7_1__20,linha7_1__19,linha7_1__18,linha7_1__17,
              linha7_1__16,linha7_1__15,linha7_1__14,linha7_1__13,linha7_1__12,
              linha7_1__11,linha7_1__10,linha7_1__9,linha7_1__8,linha7_1__7,
              linha7_1__6,linha7_1__5,linha7_1__4,linha7_1__3,linha7_1__2,
              linha7_1__1,linha7_1__0}), .a0 ({linha6_1__31,linha6_1__30,
              linha6_1__29,linha6_1__28,linha6_1__27,linha6_1__26,linha6_1__25,
              linha6_1__24,linha6_1__23,linha6_1__22,linha6_1__21,linha6_1__20,
              linha6_1__19,linha6_1__18,linha6_1__17,linha6_1__16,linha6_1__15,
              linha6_1__14,linha6_1__13,linha6_1__12,linha6_1__11,linha6_1__10,
              linha6_1__9,linha6_1__8,linha6_1__7,linha6_1__6,linha6_1__5,
              linha6_1__4,linha6_1__3,linha6_1__2,linha6_1__1,linha6_1__0}), .s (
              row_1_rowi_bni3_l)) ;
    Mux2x1_32 row_1_rowi_bni3_muxMin (.r ({linha7_2__31,linha7_2__30,
              linha7_2__29,linha7_2__28,linha7_2__27,linha7_2__26,linha7_2__25,
              linha7_2__24,linha7_2__23,linha7_2__22,linha7_2__21,linha7_2__20,
              linha7_2__19,linha7_2__18,linha7_2__17,linha7_2__16,linha7_2__15,
              linha7_2__14,linha7_2__13,linha7_2__12,linha7_2__11,linha7_2__10,
              linha7_2__9,linha7_2__8,linha7_2__7,linha7_2__6,linha7_2__5,
              linha7_2__4,linha7_2__3,linha7_2__2,linha7_2__1,linha7_2__0}), .a1 (
              {linha6_1__31,linha6_1__30,linha6_1__29,linha6_1__28,linha6_1__27,
              linha6_1__26,linha6_1__25,linha6_1__24,linha6_1__23,linha6_1__22,
              linha6_1__21,linha6_1__20,linha6_1__19,linha6_1__18,linha6_1__17,
              linha6_1__16,linha6_1__15,linha6_1__14,linha6_1__13,linha6_1__12,
              linha6_1__11,linha6_1__10,linha6_1__9,linha6_1__8,linha6_1__7,
              linha6_1__6,linha6_1__5,linha6_1__4,linha6_1__3,linha6_1__2,
              linha6_1__1,linha6_1__0}), .a0 ({linha7_1__31,linha7_1__30,
              linha7_1__29,linha7_1__28,linha7_1__27,linha7_1__26,linha7_1__25,
              linha7_1__24,linha7_1__23,linha7_1__22,linha7_1__21,linha7_1__20,
              linha7_1__19,linha7_1__18,linha7_1__17,linha7_1__16,linha7_1__15,
              linha7_1__14,linha7_1__13,linha7_1__12,linha7_1__11,linha7_1__10,
              linha7_1__9,linha7_1__8,linha7_1__7,linha7_1__6,linha7_1__5,
              linha7_1__4,linha7_1__3,linha7_1__2,linha7_1__1,linha7_1__0}), .s (
              row_1_rowi_bni3_l)) ;
    juntarComparadores_32 row_2_rowp_bni1_Comp (.g (\$dummy [7]), .l (
                          row_2_rowp_bni1_l), .a ({linha1_1__31,linha1_1__30,
                          linha1_1__29,linha1_1__28,linha1_1__27,linha1_1__26,
                          linha1_1__25,linha1_1__24,linha1_1__23,linha1_1__22,
                          linha1_1__21,linha1_1__20,linha1_1__19,linha1_1__18,
                          linha1_1__17,linha1_1__16,linha1_1__15,linha1_1__14,
                          linha1_1__13,linha1_1__12,linha1_1__11,linha1_1__10,
                          linha1_1__9,linha1_1__8,linha1_1__7,linha1_1__6,
                          linha1_1__5,linha1_1__4,linha1_1__3,linha1_1__2,
                          linha1_1__1,linha1_1__0}), .b ({linha2_2__31,
                          linha2_2__30,linha2_2__29,linha2_2__28,linha2_2__27,
                          linha2_2__26,linha2_2__25,linha2_2__24,linha2_2__23,
                          linha2_2__22,linha2_2__21,linha2_2__20,linha2_2__19,
                          linha2_2__18,linha2_2__17,linha2_2__16,linha2_2__15,
                          linha2_2__14,linha2_2__13,linha2_2__12,linha2_2__11,
                          linha2_2__10,linha2_2__9,linha2_2__8,linha2_2__7,
                          linha2_2__6,linha2_2__5,linha2_2__4,linha2_2__3,
                          linha2_2__2,linha2_2__1,linha2_2__0})) ;
    Mux2x1_32 row_2_rowp_bni1_muxMax (.r ({linha1_2__31,linha1_2__30,
              linha1_2__29,linha1_2__28,linha1_2__27,linha1_2__26,linha1_2__25,
              linha1_2__24,linha1_2__23,linha1_2__22,linha1_2__21,linha1_2__20,
              linha1_2__19,linha1_2__18,linha1_2__17,linha1_2__16,linha1_2__15,
              linha1_2__14,linha1_2__13,linha1_2__12,linha1_2__11,linha1_2__10,
              linha1_2__9,linha1_2__8,linha1_2__7,linha1_2__6,linha1_2__5,
              linha1_2__4,linha1_2__3,linha1_2__2,linha1_2__1,linha1_2__0}), .a1 (
              {linha2_2__31,linha2_2__30,linha2_2__29,linha2_2__28,linha2_2__27,
              linha2_2__26,linha2_2__25,linha2_2__24,linha2_2__23,linha2_2__22,
              linha2_2__21,linha2_2__20,linha2_2__19,linha2_2__18,linha2_2__17,
              linha2_2__16,linha2_2__15,linha2_2__14,linha2_2__13,linha2_2__12,
              linha2_2__11,linha2_2__10,linha2_2__9,linha2_2__8,linha2_2__7,
              linha2_2__6,linha2_2__5,linha2_2__4,linha2_2__3,linha2_2__2,
              linha2_2__1,linha2_2__0}), .a0 ({linha1_1__31,linha1_1__30,
              linha1_1__29,linha1_1__28,linha1_1__27,linha1_1__26,linha1_1__25,
              linha1_1__24,linha1_1__23,linha1_1__22,linha1_1__21,linha1_1__20,
              linha1_1__19,linha1_1__18,linha1_1__17,linha1_1__16,linha1_1__15,
              linha1_1__14,linha1_1__13,linha1_1__12,linha1_1__11,linha1_1__10,
              linha1_1__9,linha1_1__8,linha1_1__7,linha1_1__6,linha1_1__5,
              linha1_1__4,linha1_1__3,linha1_1__2,linha1_1__1,linha1_1__0}), .s (
              row_2_rowp_bni1_l)) ;
    Mux2x1_32 row_2_rowp_bni1_muxMin (.r ({linha2_3__31,linha2_3__30,
              linha2_3__29,linha2_3__28,linha2_3__27,linha2_3__26,linha2_3__25,
              linha2_3__24,linha2_3__23,linha2_3__22,linha2_3__21,linha2_3__20,
              linha2_3__19,linha2_3__18,linha2_3__17,linha2_3__16,linha2_3__15,
              linha2_3__14,linha2_3__13,linha2_3__12,linha2_3__11,linha2_3__10,
              linha2_3__9,linha2_3__8,linha2_3__7,linha2_3__6,linha2_3__5,
              linha2_3__4,linha2_3__3,linha2_3__2,linha2_3__1,linha2_3__0}), .a1 (
              {linha1_1__31,linha1_1__30,linha1_1__29,linha1_1__28,linha1_1__27,
              linha1_1__26,linha1_1__25,linha1_1__24,linha1_1__23,linha1_1__22,
              linha1_1__21,linha1_1__20,linha1_1__19,linha1_1__18,linha1_1__17,
              linha1_1__16,linha1_1__15,linha1_1__14,linha1_1__13,linha1_1__12,
              linha1_1__11,linha1_1__10,linha1_1__9,linha1_1__8,linha1_1__7,
              linha1_1__6,linha1_1__5,linha1_1__4,linha1_1__3,linha1_1__2,
              linha1_1__1,linha1_1__0}), .a0 ({linha2_2__31,linha2_2__30,
              linha2_2__29,linha2_2__28,linha2_2__27,linha2_2__26,linha2_2__25,
              linha2_2__24,linha2_2__23,linha2_2__22,linha2_2__21,linha2_2__20,
              linha2_2__19,linha2_2__18,linha2_2__17,linha2_2__16,linha2_2__15,
              linha2_2__14,linha2_2__13,linha2_2__12,linha2_2__11,linha2_2__10,
              linha2_2__9,linha2_2__8,linha2_2__7,linha2_2__6,linha2_2__5,
              linha2_2__4,linha2_2__3,linha2_2__2,linha2_2__1,linha2_2__0}), .s (
              row_2_rowp_bni1_l)) ;
    juntarComparadores_32 row_2_rowp_bni2_Comp (.g (\$dummy [8]), .l (
                          row_2_rowp_bni2_l), .a ({linha3_2__31,linha3_2__30,
                          linha3_2__29,linha3_2__28,linha3_2__27,linha3_2__26,
                          linha3_2__25,linha3_2__24,linha3_2__23,linha3_2__22,
                          linha3_2__21,linha3_2__20,linha3_2__19,linha3_2__18,
                          linha3_2__17,linha3_2__16,linha3_2__15,linha3_2__14,
                          linha3_2__13,linha3_2__12,linha3_2__11,linha3_2__10,
                          linha3_2__9,linha3_2__8,linha3_2__7,linha3_2__6,
                          linha3_2__5,linha3_2__4,linha3_2__3,linha3_2__2,
                          linha3_2__1,linha3_2__0}), .b ({linha4_2__31,
                          linha4_2__30,linha4_2__29,linha4_2__28,linha4_2__27,
                          linha4_2__26,linha4_2__25,linha4_2__24,linha4_2__23,
                          linha4_2__22,linha4_2__21,linha4_2__20,linha4_2__19,
                          linha4_2__18,linha4_2__17,linha4_2__16,linha4_2__15,
                          linha4_2__14,linha4_2__13,linha4_2__12,linha4_2__11,
                          linha4_2__10,linha4_2__9,linha4_2__8,linha4_2__7,
                          linha4_2__6,linha4_2__5,linha4_2__4,linha4_2__3,
                          linha4_2__2,linha4_2__1,linha4_2__0})) ;
    Mux2x1_32 row_2_rowp_bni2_muxMax (.r ({linha3_3__31,linha3_3__30,
              linha3_3__29,linha3_3__28,linha3_3__27,linha3_3__26,linha3_3__25,
              linha3_3__24,linha3_3__23,linha3_3__22,linha3_3__21,linha3_3__20,
              linha3_3__19,linha3_3__18,linha3_3__17,linha3_3__16,linha3_3__15,
              linha3_3__14,linha3_3__13,linha3_3__12,linha3_3__11,linha3_3__10,
              linha3_3__9,linha3_3__8,linha3_3__7,linha3_3__6,linha3_3__5,
              linha3_3__4,linha3_3__3,linha3_3__2,linha3_3__1,linha3_3__0}), .a1 (
              {linha4_2__31,linha4_2__30,linha4_2__29,linha4_2__28,linha4_2__27,
              linha4_2__26,linha4_2__25,linha4_2__24,linha4_2__23,linha4_2__22,
              linha4_2__21,linha4_2__20,linha4_2__19,linha4_2__18,linha4_2__17,
              linha4_2__16,linha4_2__15,linha4_2__14,linha4_2__13,linha4_2__12,
              linha4_2__11,linha4_2__10,linha4_2__9,linha4_2__8,linha4_2__7,
              linha4_2__6,linha4_2__5,linha4_2__4,linha4_2__3,linha4_2__2,
              linha4_2__1,linha4_2__0}), .a0 ({linha3_2__31,linha3_2__30,
              linha3_2__29,linha3_2__28,linha3_2__27,linha3_2__26,linha3_2__25,
              linha3_2__24,linha3_2__23,linha3_2__22,linha3_2__21,linha3_2__20,
              linha3_2__19,linha3_2__18,linha3_2__17,linha3_2__16,linha3_2__15,
              linha3_2__14,linha3_2__13,linha3_2__12,linha3_2__11,linha3_2__10,
              linha3_2__9,linha3_2__8,linha3_2__7,linha3_2__6,linha3_2__5,
              linha3_2__4,linha3_2__3,linha3_2__2,linha3_2__1,linha3_2__0}), .s (
              row_2_rowp_bni2_l)) ;
    Mux2x1_32 row_2_rowp_bni2_muxMin (.r ({linha4_3__31,linha4_3__30,
              linha4_3__29,linha4_3__28,linha4_3__27,linha4_3__26,linha4_3__25,
              linha4_3__24,linha4_3__23,linha4_3__22,linha4_3__21,linha4_3__20,
              linha4_3__19,linha4_3__18,linha4_3__17,linha4_3__16,linha4_3__15,
              linha4_3__14,linha4_3__13,linha4_3__12,linha4_3__11,linha4_3__10,
              linha4_3__9,linha4_3__8,linha4_3__7,linha4_3__6,linha4_3__5,
              linha4_3__4,linha4_3__3,linha4_3__2,linha4_3__1,linha4_3__0}), .a1 (
              {linha3_2__31,linha3_2__30,linha3_2__29,linha3_2__28,linha3_2__27,
              linha3_2__26,linha3_2__25,linha3_2__24,linha3_2__23,linha3_2__22,
              linha3_2__21,linha3_2__20,linha3_2__19,linha3_2__18,linha3_2__17,
              linha3_2__16,linha3_2__15,linha3_2__14,linha3_2__13,linha3_2__12,
              linha3_2__11,linha3_2__10,linha3_2__9,linha3_2__8,linha3_2__7,
              linha3_2__6,linha3_2__5,linha3_2__4,linha3_2__3,linha3_2__2,
              linha3_2__1,linha3_2__0}), .a0 ({linha4_2__31,linha4_2__30,
              linha4_2__29,linha4_2__28,linha4_2__27,linha4_2__26,linha4_2__25,
              linha4_2__24,linha4_2__23,linha4_2__22,linha4_2__21,linha4_2__20,
              linha4_2__19,linha4_2__18,linha4_2__17,linha4_2__16,linha4_2__15,
              linha4_2__14,linha4_2__13,linha4_2__12,linha4_2__11,linha4_2__10,
              linha4_2__9,linha4_2__8,linha4_2__7,linha4_2__6,linha4_2__5,
              linha4_2__4,linha4_2__3,linha4_2__2,linha4_2__1,linha4_2__0}), .s (
              row_2_rowp_bni2_l)) ;
    juntarComparadores_32 row_2_rowp_bni3_Comp (.g (\$dummy [9]), .l (
                          row_2_rowp_bni3_l), .a ({linha5_2__31,linha5_2__30,
                          linha5_2__29,linha5_2__28,linha5_2__27,linha5_2__26,
                          linha5_2__25,linha5_2__24,linha5_2__23,linha5_2__22,
                          linha5_2__21,linha5_2__20,linha5_2__19,linha5_2__18,
                          linha5_2__17,linha5_2__16,linha5_2__15,linha5_2__14,
                          linha5_2__13,linha5_2__12,linha5_2__11,linha5_2__10,
                          linha5_2__9,linha5_2__8,linha5_2__7,linha5_2__6,
                          linha5_2__5,linha5_2__4,linha5_2__3,linha5_2__2,
                          linha5_2__1,linha5_2__0}), .b ({linha6_2__31,
                          linha6_2__30,linha6_2__29,linha6_2__28,linha6_2__27,
                          linha6_2__26,linha6_2__25,linha6_2__24,linha6_2__23,
                          linha6_2__22,linha6_2__21,linha6_2__20,linha6_2__19,
                          linha6_2__18,linha6_2__17,linha6_2__16,linha6_2__15,
                          linha6_2__14,linha6_2__13,linha6_2__12,linha6_2__11,
                          linha6_2__10,linha6_2__9,linha6_2__8,linha6_2__7,
                          linha6_2__6,linha6_2__5,linha6_2__4,linha6_2__3,
                          linha6_2__2,linha6_2__1,linha6_2__0})) ;
    Mux2x1_32 row_2_rowp_bni3_muxMax (.r ({linha5_3__31,linha5_3__30,
              linha5_3__29,linha5_3__28,linha5_3__27,linha5_3__26,linha5_3__25,
              linha5_3__24,linha5_3__23,linha5_3__22,linha5_3__21,linha5_3__20,
              linha5_3__19,linha5_3__18,linha5_3__17,linha5_3__16,linha5_3__15,
              linha5_3__14,linha5_3__13,linha5_3__12,linha5_3__11,linha5_3__10,
              linha5_3__9,linha5_3__8,linha5_3__7,linha5_3__6,linha5_3__5,
              linha5_3__4,linha5_3__3,linha5_3__2,linha5_3__1,linha5_3__0}), .a1 (
              {linha6_2__31,linha6_2__30,linha6_2__29,linha6_2__28,linha6_2__27,
              linha6_2__26,linha6_2__25,linha6_2__24,linha6_2__23,linha6_2__22,
              linha6_2__21,linha6_2__20,linha6_2__19,linha6_2__18,linha6_2__17,
              linha6_2__16,linha6_2__15,linha6_2__14,linha6_2__13,linha6_2__12,
              linha6_2__11,linha6_2__10,linha6_2__9,linha6_2__8,linha6_2__7,
              linha6_2__6,linha6_2__5,linha6_2__4,linha6_2__3,linha6_2__2,
              linha6_2__1,linha6_2__0}), .a0 ({linha5_2__31,linha5_2__30,
              linha5_2__29,linha5_2__28,linha5_2__27,linha5_2__26,linha5_2__25,
              linha5_2__24,linha5_2__23,linha5_2__22,linha5_2__21,linha5_2__20,
              linha5_2__19,linha5_2__18,linha5_2__17,linha5_2__16,linha5_2__15,
              linha5_2__14,linha5_2__13,linha5_2__12,linha5_2__11,linha5_2__10,
              linha5_2__9,linha5_2__8,linha5_2__7,linha5_2__6,linha5_2__5,
              linha5_2__4,linha5_2__3,linha5_2__2,linha5_2__1,linha5_2__0}), .s (
              row_2_rowp_bni3_l)) ;
    Mux2x1_32 row_2_rowp_bni3_muxMin (.r ({linha6_3__31,linha6_3__30,
              linha6_3__29,linha6_3__28,linha6_3__27,linha6_3__26,linha6_3__25,
              linha6_3__24,linha6_3__23,linha6_3__22,linha6_3__21,linha6_3__20,
              linha6_3__19,linha6_3__18,linha6_3__17,linha6_3__16,linha6_3__15,
              linha6_3__14,linha6_3__13,linha6_3__12,linha6_3__11,linha6_3__10,
              linha6_3__9,linha6_3__8,linha6_3__7,linha6_3__6,linha6_3__5,
              linha6_3__4,linha6_3__3,linha6_3__2,linha6_3__1,linha6_3__0}), .a1 (
              {linha5_2__31,linha5_2__30,linha5_2__29,linha5_2__28,linha5_2__27,
              linha5_2__26,linha5_2__25,linha5_2__24,linha5_2__23,linha5_2__22,
              linha5_2__21,linha5_2__20,linha5_2__19,linha5_2__18,linha5_2__17,
              linha5_2__16,linha5_2__15,linha5_2__14,linha5_2__13,linha5_2__12,
              linha5_2__11,linha5_2__10,linha5_2__9,linha5_2__8,linha5_2__7,
              linha5_2__6,linha5_2__5,linha5_2__4,linha5_2__3,linha5_2__2,
              linha5_2__1,linha5_2__0}), .a0 ({linha6_2__31,linha6_2__30,
              linha6_2__29,linha6_2__28,linha6_2__27,linha6_2__26,linha6_2__25,
              linha6_2__24,linha6_2__23,linha6_2__22,linha6_2__21,linha6_2__20,
              linha6_2__19,linha6_2__18,linha6_2__17,linha6_2__16,linha6_2__15,
              linha6_2__14,linha6_2__13,linha6_2__12,linha6_2__11,linha6_2__10,
              linha6_2__9,linha6_2__8,linha6_2__7,linha6_2__6,linha6_2__5,
              linha6_2__4,linha6_2__3,linha6_2__2,linha6_2__1,linha6_2__0}), .s (
              row_2_rowp_bni3_l)) ;
    juntarComparadores_32 row_2_rowp_bni4_Comp (.g (\$dummy [10]), .l (
                          row_2_rowp_bni4_l), .a ({linha7_2__31,linha7_2__30,
                          linha7_2__29,linha7_2__28,linha7_2__27,linha7_2__26,
                          linha7_2__25,linha7_2__24,linha7_2__23,linha7_2__22,
                          linha7_2__21,linha7_2__20,linha7_2__19,linha7_2__18,
                          linha7_2__17,linha7_2__16,linha7_2__15,linha7_2__14,
                          linha7_2__13,linha7_2__12,linha7_2__11,linha7_2__10,
                          linha7_2__9,linha7_2__8,linha7_2__7,linha7_2__6,
                          linha7_2__5,linha7_2__4,linha7_2__3,linha7_2__2,
                          linha7_2__1,linha7_2__0}), .b ({linha8_1__31,
                          linha8_1__30,linha8_1__29,linha8_1__28,linha8_1__27,
                          linha8_1__26,linha8_1__25,linha8_1__24,linha8_1__23,
                          linha8_1__22,linha8_1__21,linha8_1__20,linha8_1__19,
                          linha8_1__18,linha8_1__17,linha8_1__16,linha8_1__15,
                          linha8_1__14,linha8_1__13,linha8_1__12,linha8_1__11,
                          linha8_1__10,linha8_1__9,linha8_1__8,linha8_1__7,
                          linha8_1__6,linha8_1__5,linha8_1__4,linha8_1__3,
                          linha8_1__2,linha8_1__1,linha8_1__0})) ;
    Mux2x1_32 row_2_rowp_bni4_muxMax (.r ({linha7_3__31,linha7_3__30,
              linha7_3__29,linha7_3__28,linha7_3__27,linha7_3__26,linha7_3__25,
              linha7_3__24,linha7_3__23,linha7_3__22,linha7_3__21,linha7_3__20,
              linha7_3__19,linha7_3__18,linha7_3__17,linha7_3__16,linha7_3__15,
              linha7_3__14,linha7_3__13,linha7_3__12,linha7_3__11,linha7_3__10,
              linha7_3__9,linha7_3__8,linha7_3__7,linha7_3__6,linha7_3__5,
              linha7_3__4,linha7_3__3,linha7_3__2,linha7_3__1,linha7_3__0}), .a1 (
              {linha8_1__31,linha8_1__30,linha8_1__29,linha8_1__28,linha8_1__27,
              linha8_1__26,linha8_1__25,linha8_1__24,linha8_1__23,linha8_1__22,
              linha8_1__21,linha8_1__20,linha8_1__19,linha8_1__18,linha8_1__17,
              linha8_1__16,linha8_1__15,linha8_1__14,linha8_1__13,linha8_1__12,
              linha8_1__11,linha8_1__10,linha8_1__9,linha8_1__8,linha8_1__7,
              linha8_1__6,linha8_1__5,linha8_1__4,linha8_1__3,linha8_1__2,
              linha8_1__1,linha8_1__0}), .a0 ({linha7_2__31,linha7_2__30,
              linha7_2__29,linha7_2__28,linha7_2__27,linha7_2__26,linha7_2__25,
              linha7_2__24,linha7_2__23,linha7_2__22,linha7_2__21,linha7_2__20,
              linha7_2__19,linha7_2__18,linha7_2__17,linha7_2__16,linha7_2__15,
              linha7_2__14,linha7_2__13,linha7_2__12,linha7_2__11,linha7_2__10,
              linha7_2__9,linha7_2__8,linha7_2__7,linha7_2__6,linha7_2__5,
              linha7_2__4,linha7_2__3,linha7_2__2,linha7_2__1,linha7_2__0}), .s (
              row_2_rowp_bni4_l)) ;
    Mux2x1_32 row_2_rowp_bni4_muxMin (.r ({linha8_2__31,linha8_2__30,
              linha8_2__29,linha8_2__28,linha8_2__27,linha8_2__26,linha8_2__25,
              linha8_2__24,linha8_2__23,linha8_2__22,linha8_2__21,linha8_2__20,
              linha8_2__19,linha8_2__18,linha8_2__17,linha8_2__16,linha8_2__15,
              linha8_2__14,linha8_2__13,linha8_2__12,linha8_2__11,linha8_2__10,
              linha8_2__9,linha8_2__8,linha8_2__7,linha8_2__6,linha8_2__5,
              linha8_2__4,linha8_2__3,linha8_2__2,linha8_2__1,linha8_2__0}), .a1 (
              {linha7_2__31,linha7_2__30,linha7_2__29,linha7_2__28,linha7_2__27,
              linha7_2__26,linha7_2__25,linha7_2__24,linha7_2__23,linha7_2__22,
              linha7_2__21,linha7_2__20,linha7_2__19,linha7_2__18,linha7_2__17,
              linha7_2__16,linha7_2__15,linha7_2__14,linha7_2__13,linha7_2__12,
              linha7_2__11,linha7_2__10,linha7_2__9,linha7_2__8,linha7_2__7,
              linha7_2__6,linha7_2__5,linha7_2__4,linha7_2__3,linha7_2__2,
              linha7_2__1,linha7_2__0}), .a0 ({linha8_1__31,linha8_1__30,
              linha8_1__29,linha8_1__28,linha8_1__27,linha8_1__26,linha8_1__25,
              linha8_1__24,linha8_1__23,linha8_1__22,linha8_1__21,linha8_1__20,
              linha8_1__19,linha8_1__18,linha8_1__17,linha8_1__16,linha8_1__15,
              linha8_1__14,linha8_1__13,linha8_1__12,linha8_1__11,linha8_1__10,
              linha8_1__9,linha8_1__8,linha8_1__7,linha8_1__6,linha8_1__5,
              linha8_1__4,linha8_1__3,linha8_1__2,linha8_1__1,linha8_1__0}), .s (
              row_2_rowp_bni4_l)) ;
    juntarComparadores_32 row_3_rowi_bni1_Comp (.g (\$dummy [11]), .l (
                          row_3_rowi_bni1_l), .a ({linha2_3__31,linha2_3__30,
                          linha2_3__29,linha2_3__28,linha2_3__27,linha2_3__26,
                          linha2_3__25,linha2_3__24,linha2_3__23,linha2_3__22,
                          linha2_3__21,linha2_3__20,linha2_3__19,linha2_3__18,
                          linha2_3__17,linha2_3__16,linha2_3__15,linha2_3__14,
                          linha2_3__13,linha2_3__12,linha2_3__11,linha2_3__10,
                          linha2_3__9,linha2_3__8,linha2_3__7,linha2_3__6,
                          linha2_3__5,linha2_3__4,linha2_3__3,linha2_3__2,
                          linha2_3__1,linha2_3__0}), .b ({linha3_3__31,
                          linha3_3__30,linha3_3__29,linha3_3__28,linha3_3__27,
                          linha3_3__26,linha3_3__25,linha3_3__24,linha3_3__23,
                          linha3_3__22,linha3_3__21,linha3_3__20,linha3_3__19,
                          linha3_3__18,linha3_3__17,linha3_3__16,linha3_3__15,
                          linha3_3__14,linha3_3__13,linha3_3__12,linha3_3__11,
                          linha3_3__10,linha3_3__9,linha3_3__8,linha3_3__7,
                          linha3_3__6,linha3_3__5,linha3_3__4,linha3_3__3,
                          linha3_3__2,linha3_3__1,linha3_3__0})) ;
    Mux2x1_32 row_3_rowi_bni1_muxMax (.r ({linha2_4__31,linha2_4__30,
              linha2_4__29,linha2_4__28,linha2_4__27,linha2_4__26,linha2_4__25,
              linha2_4__24,linha2_4__23,linha2_4__22,linha2_4__21,linha2_4__20,
              linha2_4__19,linha2_4__18,linha2_4__17,linha2_4__16,linha2_4__15,
              linha2_4__14,linha2_4__13,linha2_4__12,linha2_4__11,linha2_4__10,
              linha2_4__9,linha2_4__8,linha2_4__7,linha2_4__6,linha2_4__5,
              linha2_4__4,linha2_4__3,linha2_4__2,linha2_4__1,linha2_4__0}), .a1 (
              {linha3_3__31,linha3_3__30,linha3_3__29,linha3_3__28,linha3_3__27,
              linha3_3__26,linha3_3__25,linha3_3__24,linha3_3__23,linha3_3__22,
              linha3_3__21,linha3_3__20,linha3_3__19,linha3_3__18,linha3_3__17,
              linha3_3__16,linha3_3__15,linha3_3__14,linha3_3__13,linha3_3__12,
              linha3_3__11,linha3_3__10,linha3_3__9,linha3_3__8,linha3_3__7,
              linha3_3__6,linha3_3__5,linha3_3__4,linha3_3__3,linha3_3__2,
              linha3_3__1,linha3_3__0}), .a0 ({linha2_3__31,linha2_3__30,
              linha2_3__29,linha2_3__28,linha2_3__27,linha2_3__26,linha2_3__25,
              linha2_3__24,linha2_3__23,linha2_3__22,linha2_3__21,linha2_3__20,
              linha2_3__19,linha2_3__18,linha2_3__17,linha2_3__16,linha2_3__15,
              linha2_3__14,linha2_3__13,linha2_3__12,linha2_3__11,linha2_3__10,
              linha2_3__9,linha2_3__8,linha2_3__7,linha2_3__6,linha2_3__5,
              linha2_3__4,linha2_3__3,linha2_3__2,linha2_3__1,linha2_3__0}), .s (
              row_3_rowi_bni1_l)) ;
    Mux2x1_32 row_3_rowi_bni1_muxMin (.r ({linha3_4__31,linha3_4__30,
              linha3_4__29,linha3_4__28,linha3_4__27,linha3_4__26,linha3_4__25,
              linha3_4__24,linha3_4__23,linha3_4__22,linha3_4__21,linha3_4__20,
              linha3_4__19,linha3_4__18,linha3_4__17,linha3_4__16,linha3_4__15,
              linha3_4__14,linha3_4__13,linha3_4__12,linha3_4__11,linha3_4__10,
              linha3_4__9,linha3_4__8,linha3_4__7,linha3_4__6,linha3_4__5,
              linha3_4__4,linha3_4__3,linha3_4__2,linha3_4__1,linha3_4__0}), .a1 (
              {linha2_3__31,linha2_3__30,linha2_3__29,linha2_3__28,linha2_3__27,
              linha2_3__26,linha2_3__25,linha2_3__24,linha2_3__23,linha2_3__22,
              linha2_3__21,linha2_3__20,linha2_3__19,linha2_3__18,linha2_3__17,
              linha2_3__16,linha2_3__15,linha2_3__14,linha2_3__13,linha2_3__12,
              linha2_3__11,linha2_3__10,linha2_3__9,linha2_3__8,linha2_3__7,
              linha2_3__6,linha2_3__5,linha2_3__4,linha2_3__3,linha2_3__2,
              linha2_3__1,linha2_3__0}), .a0 ({linha3_3__31,linha3_3__30,
              linha3_3__29,linha3_3__28,linha3_3__27,linha3_3__26,linha3_3__25,
              linha3_3__24,linha3_3__23,linha3_3__22,linha3_3__21,linha3_3__20,
              linha3_3__19,linha3_3__18,linha3_3__17,linha3_3__16,linha3_3__15,
              linha3_3__14,linha3_3__13,linha3_3__12,linha3_3__11,linha3_3__10,
              linha3_3__9,linha3_3__8,linha3_3__7,linha3_3__6,linha3_3__5,
              linha3_3__4,linha3_3__3,linha3_3__2,linha3_3__1,linha3_3__0}), .s (
              row_3_rowi_bni1_l)) ;
    juntarComparadores_32 row_3_rowi_bni2_Comp (.g (\$dummy [12]), .l (
                          row_3_rowi_bni2_l), .a ({linha4_3__31,linha4_3__30,
                          linha4_3__29,linha4_3__28,linha4_3__27,linha4_3__26,
                          linha4_3__25,linha4_3__24,linha4_3__23,linha4_3__22,
                          linha4_3__21,linha4_3__20,linha4_3__19,linha4_3__18,
                          linha4_3__17,linha4_3__16,linha4_3__15,linha4_3__14,
                          linha4_3__13,linha4_3__12,linha4_3__11,linha4_3__10,
                          linha4_3__9,linha4_3__8,linha4_3__7,linha4_3__6,
                          linha4_3__5,linha4_3__4,linha4_3__3,linha4_3__2,
                          linha4_3__1,linha4_3__0}), .b ({linha5_3__31,
                          linha5_3__30,linha5_3__29,linha5_3__28,linha5_3__27,
                          linha5_3__26,linha5_3__25,linha5_3__24,linha5_3__23,
                          linha5_3__22,linha5_3__21,linha5_3__20,linha5_3__19,
                          linha5_3__18,linha5_3__17,linha5_3__16,linha5_3__15,
                          linha5_3__14,linha5_3__13,linha5_3__12,linha5_3__11,
                          linha5_3__10,linha5_3__9,linha5_3__8,linha5_3__7,
                          linha5_3__6,linha5_3__5,linha5_3__4,linha5_3__3,
                          linha5_3__2,linha5_3__1,linha5_3__0})) ;
    Mux2x1_32 row_3_rowi_bni2_muxMax (.r ({linha4_4__31,linha4_4__30,
              linha4_4__29,linha4_4__28,linha4_4__27,linha4_4__26,linha4_4__25,
              linha4_4__24,linha4_4__23,linha4_4__22,linha4_4__21,linha4_4__20,
              linha4_4__19,linha4_4__18,linha4_4__17,linha4_4__16,linha4_4__15,
              linha4_4__14,linha4_4__13,linha4_4__12,linha4_4__11,linha4_4__10,
              linha4_4__9,linha4_4__8,linha4_4__7,linha4_4__6,linha4_4__5,
              linha4_4__4,linha4_4__3,linha4_4__2,linha4_4__1,linha4_4__0}), .a1 (
              {linha5_3__31,linha5_3__30,linha5_3__29,linha5_3__28,linha5_3__27,
              linha5_3__26,linha5_3__25,linha5_3__24,linha5_3__23,linha5_3__22,
              linha5_3__21,linha5_3__20,linha5_3__19,linha5_3__18,linha5_3__17,
              linha5_3__16,linha5_3__15,linha5_3__14,linha5_3__13,linha5_3__12,
              linha5_3__11,linha5_3__10,linha5_3__9,linha5_3__8,linha5_3__7,
              linha5_3__6,linha5_3__5,linha5_3__4,linha5_3__3,linha5_3__2,
              linha5_3__1,linha5_3__0}), .a0 ({linha4_3__31,linha4_3__30,
              linha4_3__29,linha4_3__28,linha4_3__27,linha4_3__26,linha4_3__25,
              linha4_3__24,linha4_3__23,linha4_3__22,linha4_3__21,linha4_3__20,
              linha4_3__19,linha4_3__18,linha4_3__17,linha4_3__16,linha4_3__15,
              linha4_3__14,linha4_3__13,linha4_3__12,linha4_3__11,linha4_3__10,
              linha4_3__9,linha4_3__8,linha4_3__7,linha4_3__6,linha4_3__5,
              linha4_3__4,linha4_3__3,linha4_3__2,linha4_3__1,linha4_3__0}), .s (
              row_3_rowi_bni2_l)) ;
    Mux2x1_32 row_3_rowi_bni2_muxMin (.r ({linha5_4__31,linha5_4__30,
              linha5_4__29,linha5_4__28,linha5_4__27,linha5_4__26,linha5_4__25,
              linha5_4__24,linha5_4__23,linha5_4__22,linha5_4__21,linha5_4__20,
              linha5_4__19,linha5_4__18,linha5_4__17,linha5_4__16,linha5_4__15,
              linha5_4__14,linha5_4__13,linha5_4__12,linha5_4__11,linha5_4__10,
              linha5_4__9,linha5_4__8,linha5_4__7,linha5_4__6,linha5_4__5,
              linha5_4__4,linha5_4__3,linha5_4__2,linha5_4__1,linha5_4__0}), .a1 (
              {linha4_3__31,linha4_3__30,linha4_3__29,linha4_3__28,linha4_3__27,
              linha4_3__26,linha4_3__25,linha4_3__24,linha4_3__23,linha4_3__22,
              linha4_3__21,linha4_3__20,linha4_3__19,linha4_3__18,linha4_3__17,
              linha4_3__16,linha4_3__15,linha4_3__14,linha4_3__13,linha4_3__12,
              linha4_3__11,linha4_3__10,linha4_3__9,linha4_3__8,linha4_3__7,
              linha4_3__6,linha4_3__5,linha4_3__4,linha4_3__3,linha4_3__2,
              linha4_3__1,linha4_3__0}), .a0 ({linha5_3__31,linha5_3__30,
              linha5_3__29,linha5_3__28,linha5_3__27,linha5_3__26,linha5_3__25,
              linha5_3__24,linha5_3__23,linha5_3__22,linha5_3__21,linha5_3__20,
              linha5_3__19,linha5_3__18,linha5_3__17,linha5_3__16,linha5_3__15,
              linha5_3__14,linha5_3__13,linha5_3__12,linha5_3__11,linha5_3__10,
              linha5_3__9,linha5_3__8,linha5_3__7,linha5_3__6,linha5_3__5,
              linha5_3__4,linha5_3__3,linha5_3__2,linha5_3__1,linha5_3__0}), .s (
              row_3_rowi_bni2_l)) ;
    juntarComparadores_32 row_3_rowi_bni3_Comp (.g (\$dummy [13]), .l (
                          row_3_rowi_bni3_l), .a ({linha6_3__31,linha6_3__30,
                          linha6_3__29,linha6_3__28,linha6_3__27,linha6_3__26,
                          linha6_3__25,linha6_3__24,linha6_3__23,linha6_3__22,
                          linha6_3__21,linha6_3__20,linha6_3__19,linha6_3__18,
                          linha6_3__17,linha6_3__16,linha6_3__15,linha6_3__14,
                          linha6_3__13,linha6_3__12,linha6_3__11,linha6_3__10,
                          linha6_3__9,linha6_3__8,linha6_3__7,linha6_3__6,
                          linha6_3__5,linha6_3__4,linha6_3__3,linha6_3__2,
                          linha6_3__1,linha6_3__0}), .b ({linha7_3__31,
                          linha7_3__30,linha7_3__29,linha7_3__28,linha7_3__27,
                          linha7_3__26,linha7_3__25,linha7_3__24,linha7_3__23,
                          linha7_3__22,linha7_3__21,linha7_3__20,linha7_3__19,
                          linha7_3__18,linha7_3__17,linha7_3__16,linha7_3__15,
                          linha7_3__14,linha7_3__13,linha7_3__12,linha7_3__11,
                          linha7_3__10,linha7_3__9,linha7_3__8,linha7_3__7,
                          linha7_3__6,linha7_3__5,linha7_3__4,linha7_3__3,
                          linha7_3__2,linha7_3__1,linha7_3__0})) ;
    Mux2x1_32 row_3_rowi_bni3_muxMax (.r ({linha6_4__31,linha6_4__30,
              linha6_4__29,linha6_4__28,linha6_4__27,linha6_4__26,linha6_4__25,
              linha6_4__24,linha6_4__23,linha6_4__22,linha6_4__21,linha6_4__20,
              linha6_4__19,linha6_4__18,linha6_4__17,linha6_4__16,linha6_4__15,
              linha6_4__14,linha6_4__13,linha6_4__12,linha6_4__11,linha6_4__10,
              linha6_4__9,linha6_4__8,linha6_4__7,linha6_4__6,linha6_4__5,
              linha6_4__4,linha6_4__3,linha6_4__2,linha6_4__1,linha6_4__0}), .a1 (
              {linha7_3__31,linha7_3__30,linha7_3__29,linha7_3__28,linha7_3__27,
              linha7_3__26,linha7_3__25,linha7_3__24,linha7_3__23,linha7_3__22,
              linha7_3__21,linha7_3__20,linha7_3__19,linha7_3__18,linha7_3__17,
              linha7_3__16,linha7_3__15,linha7_3__14,linha7_3__13,linha7_3__12,
              linha7_3__11,linha7_3__10,linha7_3__9,linha7_3__8,linha7_3__7,
              linha7_3__6,linha7_3__5,linha7_3__4,linha7_3__3,linha7_3__2,
              linha7_3__1,linha7_3__0}), .a0 ({linha6_3__31,linha6_3__30,
              linha6_3__29,linha6_3__28,linha6_3__27,linha6_3__26,linha6_3__25,
              linha6_3__24,linha6_3__23,linha6_3__22,linha6_3__21,linha6_3__20,
              linha6_3__19,linha6_3__18,linha6_3__17,linha6_3__16,linha6_3__15,
              linha6_3__14,linha6_3__13,linha6_3__12,linha6_3__11,linha6_3__10,
              linha6_3__9,linha6_3__8,linha6_3__7,linha6_3__6,linha6_3__5,
              linha6_3__4,linha6_3__3,linha6_3__2,linha6_3__1,linha6_3__0}), .s (
              row_3_rowi_bni3_l)) ;
    Mux2x1_32 row_3_rowi_bni3_muxMin (.r ({linha7_4__31,linha7_4__30,
              linha7_4__29,linha7_4__28,linha7_4__27,linha7_4__26,linha7_4__25,
              linha7_4__24,linha7_4__23,linha7_4__22,linha7_4__21,linha7_4__20,
              linha7_4__19,linha7_4__18,linha7_4__17,linha7_4__16,linha7_4__15,
              linha7_4__14,linha7_4__13,linha7_4__12,linha7_4__11,linha7_4__10,
              linha7_4__9,linha7_4__8,linha7_4__7,linha7_4__6,linha7_4__5,
              linha7_4__4,linha7_4__3,linha7_4__2,linha7_4__1,linha7_4__0}), .a1 (
              {linha6_3__31,linha6_3__30,linha6_3__29,linha6_3__28,linha6_3__27,
              linha6_3__26,linha6_3__25,linha6_3__24,linha6_3__23,linha6_3__22,
              linha6_3__21,linha6_3__20,linha6_3__19,linha6_3__18,linha6_3__17,
              linha6_3__16,linha6_3__15,linha6_3__14,linha6_3__13,linha6_3__12,
              linha6_3__11,linha6_3__10,linha6_3__9,linha6_3__8,linha6_3__7,
              linha6_3__6,linha6_3__5,linha6_3__4,linha6_3__3,linha6_3__2,
              linha6_3__1,linha6_3__0}), .a0 ({linha7_3__31,linha7_3__30,
              linha7_3__29,linha7_3__28,linha7_3__27,linha7_3__26,linha7_3__25,
              linha7_3__24,linha7_3__23,linha7_3__22,linha7_3__21,linha7_3__20,
              linha7_3__19,linha7_3__18,linha7_3__17,linha7_3__16,linha7_3__15,
              linha7_3__14,linha7_3__13,linha7_3__12,linha7_3__11,linha7_3__10,
              linha7_3__9,linha7_3__8,linha7_3__7,linha7_3__6,linha7_3__5,
              linha7_3__4,linha7_3__3,linha7_3__2,linha7_3__1,linha7_3__0}), .s (
              row_3_rowi_bni3_l)) ;
    juntarComparadores_32 row_4_rowp_bni1_Comp (.g (\$dummy [14]), .l (
                          row_4_rowp_bni1_l), .a ({linha1_2__31,linha1_2__30,
                          linha1_2__29,linha1_2__28,linha1_2__27,linha1_2__26,
                          linha1_2__25,linha1_2__24,linha1_2__23,linha1_2__22,
                          linha1_2__21,linha1_2__20,linha1_2__19,linha1_2__18,
                          linha1_2__17,linha1_2__16,linha1_2__15,linha1_2__14,
                          linha1_2__13,linha1_2__12,linha1_2__11,linha1_2__10,
                          linha1_2__9,linha1_2__8,linha1_2__7,linha1_2__6,
                          linha1_2__5,linha1_2__4,linha1_2__3,linha1_2__2,
                          linha1_2__1,linha1_2__0}), .b ({linha2_4__31,
                          linha2_4__30,linha2_4__29,linha2_4__28,linha2_4__27,
                          linha2_4__26,linha2_4__25,linha2_4__24,linha2_4__23,
                          linha2_4__22,linha2_4__21,linha2_4__20,linha2_4__19,
                          linha2_4__18,linha2_4__17,linha2_4__16,linha2_4__15,
                          linha2_4__14,linha2_4__13,linha2_4__12,linha2_4__11,
                          linha2_4__10,linha2_4__9,linha2_4__8,linha2_4__7,
                          linha2_4__6,linha2_4__5,linha2_4__4,linha2_4__3,
                          linha2_4__2,linha2_4__1,linha2_4__0})) ;
    Mux2x1_32 row_4_rowp_bni1_muxMax (.r ({linha1_3__31,linha1_3__30,
              linha1_3__29,linha1_3__28,linha1_3__27,linha1_3__26,linha1_3__25,
              linha1_3__24,linha1_3__23,linha1_3__22,linha1_3__21,linha1_3__20,
              linha1_3__19,linha1_3__18,linha1_3__17,linha1_3__16,linha1_3__15,
              linha1_3__14,linha1_3__13,linha1_3__12,linha1_3__11,linha1_3__10,
              linha1_3__9,linha1_3__8,linha1_3__7,linha1_3__6,linha1_3__5,
              linha1_3__4,linha1_3__3,linha1_3__2,linha1_3__1,linha1_3__0}), .a1 (
              {linha2_4__31,linha2_4__30,linha2_4__29,linha2_4__28,linha2_4__27,
              linha2_4__26,linha2_4__25,linha2_4__24,linha2_4__23,linha2_4__22,
              linha2_4__21,linha2_4__20,linha2_4__19,linha2_4__18,linha2_4__17,
              linha2_4__16,linha2_4__15,linha2_4__14,linha2_4__13,linha2_4__12,
              linha2_4__11,linha2_4__10,linha2_4__9,linha2_4__8,linha2_4__7,
              linha2_4__6,linha2_4__5,linha2_4__4,linha2_4__3,linha2_4__2,
              linha2_4__1,linha2_4__0}), .a0 ({linha1_2__31,linha1_2__30,
              linha1_2__29,linha1_2__28,linha1_2__27,linha1_2__26,linha1_2__25,
              linha1_2__24,linha1_2__23,linha1_2__22,linha1_2__21,linha1_2__20,
              linha1_2__19,linha1_2__18,linha1_2__17,linha1_2__16,linha1_2__15,
              linha1_2__14,linha1_2__13,linha1_2__12,linha1_2__11,linha1_2__10,
              linha1_2__9,linha1_2__8,linha1_2__7,linha1_2__6,linha1_2__5,
              linha1_2__4,linha1_2__3,linha1_2__2,linha1_2__1,linha1_2__0}), .s (
              row_4_rowp_bni1_l)) ;
    Mux2x1_32 row_4_rowp_bni1_muxMin (.r ({linha2_5__31,linha2_5__30,
              linha2_5__29,linha2_5__28,linha2_5__27,linha2_5__26,linha2_5__25,
              linha2_5__24,linha2_5__23,linha2_5__22,linha2_5__21,linha2_5__20,
              linha2_5__19,linha2_5__18,linha2_5__17,linha2_5__16,linha2_5__15,
              linha2_5__14,linha2_5__13,linha2_5__12,linha2_5__11,linha2_5__10,
              linha2_5__9,linha2_5__8,linha2_5__7,linha2_5__6,linha2_5__5,
              linha2_5__4,linha2_5__3,linha2_5__2,linha2_5__1,linha2_5__0}), .a1 (
              {linha1_2__31,linha1_2__30,linha1_2__29,linha1_2__28,linha1_2__27,
              linha1_2__26,linha1_2__25,linha1_2__24,linha1_2__23,linha1_2__22,
              linha1_2__21,linha1_2__20,linha1_2__19,linha1_2__18,linha1_2__17,
              linha1_2__16,linha1_2__15,linha1_2__14,linha1_2__13,linha1_2__12,
              linha1_2__11,linha1_2__10,linha1_2__9,linha1_2__8,linha1_2__7,
              linha1_2__6,linha1_2__5,linha1_2__4,linha1_2__3,linha1_2__2,
              linha1_2__1,linha1_2__0}), .a0 ({linha2_4__31,linha2_4__30,
              linha2_4__29,linha2_4__28,linha2_4__27,linha2_4__26,linha2_4__25,
              linha2_4__24,linha2_4__23,linha2_4__22,linha2_4__21,linha2_4__20,
              linha2_4__19,linha2_4__18,linha2_4__17,linha2_4__16,linha2_4__15,
              linha2_4__14,linha2_4__13,linha2_4__12,linha2_4__11,linha2_4__10,
              linha2_4__9,linha2_4__8,linha2_4__7,linha2_4__6,linha2_4__5,
              linha2_4__4,linha2_4__3,linha2_4__2,linha2_4__1,linha2_4__0}), .s (
              row_4_rowp_bni1_l)) ;
    juntarComparadores_32 row_4_rowp_bni2_Comp (.g (\$dummy [15]), .l (
                          row_4_rowp_bni2_l), .a ({linha3_4__31,linha3_4__30,
                          linha3_4__29,linha3_4__28,linha3_4__27,linha3_4__26,
                          linha3_4__25,linha3_4__24,linha3_4__23,linha3_4__22,
                          linha3_4__21,linha3_4__20,linha3_4__19,linha3_4__18,
                          linha3_4__17,linha3_4__16,linha3_4__15,linha3_4__14,
                          linha3_4__13,linha3_4__12,linha3_4__11,linha3_4__10,
                          linha3_4__9,linha3_4__8,linha3_4__7,linha3_4__6,
                          linha3_4__5,linha3_4__4,linha3_4__3,linha3_4__2,
                          linha3_4__1,linha3_4__0}), .b ({linha4_4__31,
                          linha4_4__30,linha4_4__29,linha4_4__28,linha4_4__27,
                          linha4_4__26,linha4_4__25,linha4_4__24,linha4_4__23,
                          linha4_4__22,linha4_4__21,linha4_4__20,linha4_4__19,
                          linha4_4__18,linha4_4__17,linha4_4__16,linha4_4__15,
                          linha4_4__14,linha4_4__13,linha4_4__12,linha4_4__11,
                          linha4_4__10,linha4_4__9,linha4_4__8,linha4_4__7,
                          linha4_4__6,linha4_4__5,linha4_4__4,linha4_4__3,
                          linha4_4__2,linha4_4__1,linha4_4__0})) ;
    Mux2x1_32 row_4_rowp_bni2_muxMax (.r ({linha3_5__31,linha3_5__30,
              linha3_5__29,linha3_5__28,linha3_5__27,linha3_5__26,linha3_5__25,
              linha3_5__24,linha3_5__23,linha3_5__22,linha3_5__21,linha3_5__20,
              linha3_5__19,linha3_5__18,linha3_5__17,linha3_5__16,linha3_5__15,
              linha3_5__14,linha3_5__13,linha3_5__12,linha3_5__11,linha3_5__10,
              linha3_5__9,linha3_5__8,linha3_5__7,linha3_5__6,linha3_5__5,
              linha3_5__4,linha3_5__3,linha3_5__2,linha3_5__1,linha3_5__0}), .a1 (
              {linha4_4__31,linha4_4__30,linha4_4__29,linha4_4__28,linha4_4__27,
              linha4_4__26,linha4_4__25,linha4_4__24,linha4_4__23,linha4_4__22,
              linha4_4__21,linha4_4__20,linha4_4__19,linha4_4__18,linha4_4__17,
              linha4_4__16,linha4_4__15,linha4_4__14,linha4_4__13,linha4_4__12,
              linha4_4__11,linha4_4__10,linha4_4__9,linha4_4__8,linha4_4__7,
              linha4_4__6,linha4_4__5,linha4_4__4,linha4_4__3,linha4_4__2,
              linha4_4__1,linha4_4__0}), .a0 ({linha3_4__31,linha3_4__30,
              linha3_4__29,linha3_4__28,linha3_4__27,linha3_4__26,linha3_4__25,
              linha3_4__24,linha3_4__23,linha3_4__22,linha3_4__21,linha3_4__20,
              linha3_4__19,linha3_4__18,linha3_4__17,linha3_4__16,linha3_4__15,
              linha3_4__14,linha3_4__13,linha3_4__12,linha3_4__11,linha3_4__10,
              linha3_4__9,linha3_4__8,linha3_4__7,linha3_4__6,linha3_4__5,
              linha3_4__4,linha3_4__3,linha3_4__2,linha3_4__1,linha3_4__0}), .s (
              row_4_rowp_bni2_l)) ;
    Mux2x1_32 row_4_rowp_bni2_muxMin (.r ({linha4_5__31,linha4_5__30,
              linha4_5__29,linha4_5__28,linha4_5__27,linha4_5__26,linha4_5__25,
              linha4_5__24,linha4_5__23,linha4_5__22,linha4_5__21,linha4_5__20,
              linha4_5__19,linha4_5__18,linha4_5__17,linha4_5__16,linha4_5__15,
              linha4_5__14,linha4_5__13,linha4_5__12,linha4_5__11,linha4_5__10,
              linha4_5__9,linha4_5__8,linha4_5__7,linha4_5__6,linha4_5__5,
              linha4_5__4,linha4_5__3,linha4_5__2,linha4_5__1,linha4_5__0}), .a1 (
              {linha3_4__31,linha3_4__30,linha3_4__29,linha3_4__28,linha3_4__27,
              linha3_4__26,linha3_4__25,linha3_4__24,linha3_4__23,linha3_4__22,
              linha3_4__21,linha3_4__20,linha3_4__19,linha3_4__18,linha3_4__17,
              linha3_4__16,linha3_4__15,linha3_4__14,linha3_4__13,linha3_4__12,
              linha3_4__11,linha3_4__10,linha3_4__9,linha3_4__8,linha3_4__7,
              linha3_4__6,linha3_4__5,linha3_4__4,linha3_4__3,linha3_4__2,
              linha3_4__1,linha3_4__0}), .a0 ({linha4_4__31,linha4_4__30,
              linha4_4__29,linha4_4__28,linha4_4__27,linha4_4__26,linha4_4__25,
              linha4_4__24,linha4_4__23,linha4_4__22,linha4_4__21,linha4_4__20,
              linha4_4__19,linha4_4__18,linha4_4__17,linha4_4__16,linha4_4__15,
              linha4_4__14,linha4_4__13,linha4_4__12,linha4_4__11,linha4_4__10,
              linha4_4__9,linha4_4__8,linha4_4__7,linha4_4__6,linha4_4__5,
              linha4_4__4,linha4_4__3,linha4_4__2,linha4_4__1,linha4_4__0}), .s (
              row_4_rowp_bni2_l)) ;
    juntarComparadores_32 row_4_rowp_bni3_Comp (.g (\$dummy [16]), .l (
                          row_4_rowp_bni3_l), .a ({linha5_4__31,linha5_4__30,
                          linha5_4__29,linha5_4__28,linha5_4__27,linha5_4__26,
                          linha5_4__25,linha5_4__24,linha5_4__23,linha5_4__22,
                          linha5_4__21,linha5_4__20,linha5_4__19,linha5_4__18,
                          linha5_4__17,linha5_4__16,linha5_4__15,linha5_4__14,
                          linha5_4__13,linha5_4__12,linha5_4__11,linha5_4__10,
                          linha5_4__9,linha5_4__8,linha5_4__7,linha5_4__6,
                          linha5_4__5,linha5_4__4,linha5_4__3,linha5_4__2,
                          linha5_4__1,linha5_4__0}), .b ({linha6_4__31,
                          linha6_4__30,linha6_4__29,linha6_4__28,linha6_4__27,
                          linha6_4__26,linha6_4__25,linha6_4__24,linha6_4__23,
                          linha6_4__22,linha6_4__21,linha6_4__20,linha6_4__19,
                          linha6_4__18,linha6_4__17,linha6_4__16,linha6_4__15,
                          linha6_4__14,linha6_4__13,linha6_4__12,linha6_4__11,
                          linha6_4__10,linha6_4__9,linha6_4__8,linha6_4__7,
                          linha6_4__6,linha6_4__5,linha6_4__4,linha6_4__3,
                          linha6_4__2,linha6_4__1,linha6_4__0})) ;
    Mux2x1_32 row_4_rowp_bni3_muxMax (.r ({linha5_5__31,linha5_5__30,
              linha5_5__29,linha5_5__28,linha5_5__27,linha5_5__26,linha5_5__25,
              linha5_5__24,linha5_5__23,linha5_5__22,linha5_5__21,linha5_5__20,
              linha5_5__19,linha5_5__18,linha5_5__17,linha5_5__16,linha5_5__15,
              linha5_5__14,linha5_5__13,linha5_5__12,linha5_5__11,linha5_5__10,
              linha5_5__9,linha5_5__8,linha5_5__7,linha5_5__6,linha5_5__5,
              linha5_5__4,linha5_5__3,linha5_5__2,linha5_5__1,linha5_5__0}), .a1 (
              {linha6_4__31,linha6_4__30,linha6_4__29,linha6_4__28,linha6_4__27,
              linha6_4__26,linha6_4__25,linha6_4__24,linha6_4__23,linha6_4__22,
              linha6_4__21,linha6_4__20,linha6_4__19,linha6_4__18,linha6_4__17,
              linha6_4__16,linha6_4__15,linha6_4__14,linha6_4__13,linha6_4__12,
              linha6_4__11,linha6_4__10,linha6_4__9,linha6_4__8,linha6_4__7,
              linha6_4__6,linha6_4__5,linha6_4__4,linha6_4__3,linha6_4__2,
              linha6_4__1,linha6_4__0}), .a0 ({linha5_4__31,linha5_4__30,
              linha5_4__29,linha5_4__28,linha5_4__27,linha5_4__26,linha5_4__25,
              linha5_4__24,linha5_4__23,linha5_4__22,linha5_4__21,linha5_4__20,
              linha5_4__19,linha5_4__18,linha5_4__17,linha5_4__16,linha5_4__15,
              linha5_4__14,linha5_4__13,linha5_4__12,linha5_4__11,linha5_4__10,
              linha5_4__9,linha5_4__8,linha5_4__7,linha5_4__6,linha5_4__5,
              linha5_4__4,linha5_4__3,linha5_4__2,linha5_4__1,linha5_4__0}), .s (
              row_4_rowp_bni3_l)) ;
    Mux2x1_32 row_4_rowp_bni3_muxMin (.r ({linha6_5__31,linha6_5__30,
              linha6_5__29,linha6_5__28,linha6_5__27,linha6_5__26,linha6_5__25,
              linha6_5__24,linha6_5__23,linha6_5__22,linha6_5__21,linha6_5__20,
              linha6_5__19,linha6_5__18,linha6_5__17,linha6_5__16,linha6_5__15,
              linha6_5__14,linha6_5__13,linha6_5__12,linha6_5__11,linha6_5__10,
              linha6_5__9,linha6_5__8,linha6_5__7,linha6_5__6,linha6_5__5,
              linha6_5__4,linha6_5__3,linha6_5__2,linha6_5__1,linha6_5__0}), .a1 (
              {linha5_4__31,linha5_4__30,linha5_4__29,linha5_4__28,linha5_4__27,
              linha5_4__26,linha5_4__25,linha5_4__24,linha5_4__23,linha5_4__22,
              linha5_4__21,linha5_4__20,linha5_4__19,linha5_4__18,linha5_4__17,
              linha5_4__16,linha5_4__15,linha5_4__14,linha5_4__13,linha5_4__12,
              linha5_4__11,linha5_4__10,linha5_4__9,linha5_4__8,linha5_4__7,
              linha5_4__6,linha5_4__5,linha5_4__4,linha5_4__3,linha5_4__2,
              linha5_4__1,linha5_4__0}), .a0 ({linha6_4__31,linha6_4__30,
              linha6_4__29,linha6_4__28,linha6_4__27,linha6_4__26,linha6_4__25,
              linha6_4__24,linha6_4__23,linha6_4__22,linha6_4__21,linha6_4__20,
              linha6_4__19,linha6_4__18,linha6_4__17,linha6_4__16,linha6_4__15,
              linha6_4__14,linha6_4__13,linha6_4__12,linha6_4__11,linha6_4__10,
              linha6_4__9,linha6_4__8,linha6_4__7,linha6_4__6,linha6_4__5,
              linha6_4__4,linha6_4__3,linha6_4__2,linha6_4__1,linha6_4__0}), .s (
              row_4_rowp_bni3_l)) ;
    juntarComparadores_32 row_4_rowp_bni4_Comp (.g (\$dummy [17]), .l (
                          row_4_rowp_bni4_l), .a ({linha7_4__31,linha7_4__30,
                          linha7_4__29,linha7_4__28,linha7_4__27,linha7_4__26,
                          linha7_4__25,linha7_4__24,linha7_4__23,linha7_4__22,
                          linha7_4__21,linha7_4__20,linha7_4__19,linha7_4__18,
                          linha7_4__17,linha7_4__16,linha7_4__15,linha7_4__14,
                          linha7_4__13,linha7_4__12,linha7_4__11,linha7_4__10,
                          linha7_4__9,linha7_4__8,linha7_4__7,linha7_4__6,
                          linha7_4__5,linha7_4__4,linha7_4__3,linha7_4__2,
                          linha7_4__1,linha7_4__0}), .b ({linha8_2__31,
                          linha8_2__30,linha8_2__29,linha8_2__28,linha8_2__27,
                          linha8_2__26,linha8_2__25,linha8_2__24,linha8_2__23,
                          linha8_2__22,linha8_2__21,linha8_2__20,linha8_2__19,
                          linha8_2__18,linha8_2__17,linha8_2__16,linha8_2__15,
                          linha8_2__14,linha8_2__13,linha8_2__12,linha8_2__11,
                          linha8_2__10,linha8_2__9,linha8_2__8,linha8_2__7,
                          linha8_2__6,linha8_2__5,linha8_2__4,linha8_2__3,
                          linha8_2__2,linha8_2__1,linha8_2__0})) ;
    Mux2x1_32 row_4_rowp_bni4_muxMax (.r ({linha7_5__31,linha7_5__30,
              linha7_5__29,linha7_5__28,linha7_5__27,linha7_5__26,linha7_5__25,
              linha7_5__24,linha7_5__23,linha7_5__22,linha7_5__21,linha7_5__20,
              linha7_5__19,linha7_5__18,linha7_5__17,linha7_5__16,linha7_5__15,
              linha7_5__14,linha7_5__13,linha7_5__12,linha7_5__11,linha7_5__10,
              linha7_5__9,linha7_5__8,linha7_5__7,linha7_5__6,linha7_5__5,
              linha7_5__4,linha7_5__3,linha7_5__2,linha7_5__1,linha7_5__0}), .a1 (
              {linha8_2__31,linha8_2__30,linha8_2__29,linha8_2__28,linha8_2__27,
              linha8_2__26,linha8_2__25,linha8_2__24,linha8_2__23,linha8_2__22,
              linha8_2__21,linha8_2__20,linha8_2__19,linha8_2__18,linha8_2__17,
              linha8_2__16,linha8_2__15,linha8_2__14,linha8_2__13,linha8_2__12,
              linha8_2__11,linha8_2__10,linha8_2__9,linha8_2__8,linha8_2__7,
              linha8_2__6,linha8_2__5,linha8_2__4,linha8_2__3,linha8_2__2,
              linha8_2__1,linha8_2__0}), .a0 ({linha7_4__31,linha7_4__30,
              linha7_4__29,linha7_4__28,linha7_4__27,linha7_4__26,linha7_4__25,
              linha7_4__24,linha7_4__23,linha7_4__22,linha7_4__21,linha7_4__20,
              linha7_4__19,linha7_4__18,linha7_4__17,linha7_4__16,linha7_4__15,
              linha7_4__14,linha7_4__13,linha7_4__12,linha7_4__11,linha7_4__10,
              linha7_4__9,linha7_4__8,linha7_4__7,linha7_4__6,linha7_4__5,
              linha7_4__4,linha7_4__3,linha7_4__2,linha7_4__1,linha7_4__0}), .s (
              row_4_rowp_bni4_l)) ;
    Mux2x1_32 row_4_rowp_bni4_muxMin (.r ({linha8_3__31,linha8_3__30,
              linha8_3__29,linha8_3__28,linha8_3__27,linha8_3__26,linha8_3__25,
              linha8_3__24,linha8_3__23,linha8_3__22,linha8_3__21,linha8_3__20,
              linha8_3__19,linha8_3__18,linha8_3__17,linha8_3__16,linha8_3__15,
              linha8_3__14,linha8_3__13,linha8_3__12,linha8_3__11,linha8_3__10,
              linha8_3__9,linha8_3__8,linha8_3__7,linha8_3__6,linha8_3__5,
              linha8_3__4,linha8_3__3,linha8_3__2,linha8_3__1,linha8_3__0}), .a1 (
              {linha7_4__31,linha7_4__30,linha7_4__29,linha7_4__28,linha7_4__27,
              linha7_4__26,linha7_4__25,linha7_4__24,linha7_4__23,linha7_4__22,
              linha7_4__21,linha7_4__20,linha7_4__19,linha7_4__18,linha7_4__17,
              linha7_4__16,linha7_4__15,linha7_4__14,linha7_4__13,linha7_4__12,
              linha7_4__11,linha7_4__10,linha7_4__9,linha7_4__8,linha7_4__7,
              linha7_4__6,linha7_4__5,linha7_4__4,linha7_4__3,linha7_4__2,
              linha7_4__1,linha7_4__0}), .a0 ({linha8_2__31,linha8_2__30,
              linha8_2__29,linha8_2__28,linha8_2__27,linha8_2__26,linha8_2__25,
              linha8_2__24,linha8_2__23,linha8_2__22,linha8_2__21,linha8_2__20,
              linha8_2__19,linha8_2__18,linha8_2__17,linha8_2__16,linha8_2__15,
              linha8_2__14,linha8_2__13,linha8_2__12,linha8_2__11,linha8_2__10,
              linha8_2__9,linha8_2__8,linha8_2__7,linha8_2__6,linha8_2__5,
              linha8_2__4,linha8_2__3,linha8_2__2,linha8_2__1,linha8_2__0}), .s (
              row_4_rowp_bni4_l)) ;
    juntarComparadores_32 row_5_rowi_bni1_Comp (.g (\$dummy [18]), .l (
                          row_5_rowi_bni1_l), .a ({linha2_5__31,linha2_5__30,
                          linha2_5__29,linha2_5__28,linha2_5__27,linha2_5__26,
                          linha2_5__25,linha2_5__24,linha2_5__23,linha2_5__22,
                          linha2_5__21,linha2_5__20,linha2_5__19,linha2_5__18,
                          linha2_5__17,linha2_5__16,linha2_5__15,linha2_5__14,
                          linha2_5__13,linha2_5__12,linha2_5__11,linha2_5__10,
                          linha2_5__9,linha2_5__8,linha2_5__7,linha2_5__6,
                          linha2_5__5,linha2_5__4,linha2_5__3,linha2_5__2,
                          linha2_5__1,linha2_5__0}), .b ({linha3_5__31,
                          linha3_5__30,linha3_5__29,linha3_5__28,linha3_5__27,
                          linha3_5__26,linha3_5__25,linha3_5__24,linha3_5__23,
                          linha3_5__22,linha3_5__21,linha3_5__20,linha3_5__19,
                          linha3_5__18,linha3_5__17,linha3_5__16,linha3_5__15,
                          linha3_5__14,linha3_5__13,linha3_5__12,linha3_5__11,
                          linha3_5__10,linha3_5__9,linha3_5__8,linha3_5__7,
                          linha3_5__6,linha3_5__5,linha3_5__4,linha3_5__3,
                          linha3_5__2,linha3_5__1,linha3_5__0})) ;
    Mux2x1_32 row_5_rowi_bni1_muxMax (.r ({linha2_6__31,linha2_6__30,
              linha2_6__29,linha2_6__28,linha2_6__27,linha2_6__26,linha2_6__25,
              linha2_6__24,linha2_6__23,linha2_6__22,linha2_6__21,linha2_6__20,
              linha2_6__19,linha2_6__18,linha2_6__17,linha2_6__16,linha2_6__15,
              linha2_6__14,linha2_6__13,linha2_6__12,linha2_6__11,linha2_6__10,
              linha2_6__9,linha2_6__8,linha2_6__7,linha2_6__6,linha2_6__5,
              linha2_6__4,linha2_6__3,linha2_6__2,linha2_6__1,linha2_6__0}), .a1 (
              {linha3_5__31,linha3_5__30,linha3_5__29,linha3_5__28,linha3_5__27,
              linha3_5__26,linha3_5__25,linha3_5__24,linha3_5__23,linha3_5__22,
              linha3_5__21,linha3_5__20,linha3_5__19,linha3_5__18,linha3_5__17,
              linha3_5__16,linha3_5__15,linha3_5__14,linha3_5__13,linha3_5__12,
              linha3_5__11,linha3_5__10,linha3_5__9,linha3_5__8,linha3_5__7,
              linha3_5__6,linha3_5__5,linha3_5__4,linha3_5__3,linha3_5__2,
              linha3_5__1,linha3_5__0}), .a0 ({linha2_5__31,linha2_5__30,
              linha2_5__29,linha2_5__28,linha2_5__27,linha2_5__26,linha2_5__25,
              linha2_5__24,linha2_5__23,linha2_5__22,linha2_5__21,linha2_5__20,
              linha2_5__19,linha2_5__18,linha2_5__17,linha2_5__16,linha2_5__15,
              linha2_5__14,linha2_5__13,linha2_5__12,linha2_5__11,linha2_5__10,
              linha2_5__9,linha2_5__8,linha2_5__7,linha2_5__6,linha2_5__5,
              linha2_5__4,linha2_5__3,linha2_5__2,linha2_5__1,linha2_5__0}), .s (
              row_5_rowi_bni1_l)) ;
    Mux2x1_32 row_5_rowi_bni1_muxMin (.r ({linha3_6__31,linha3_6__30,
              linha3_6__29,linha3_6__28,linha3_6__27,linha3_6__26,linha3_6__25,
              linha3_6__24,linha3_6__23,linha3_6__22,linha3_6__21,linha3_6__20,
              linha3_6__19,linha3_6__18,linha3_6__17,linha3_6__16,linha3_6__15,
              linha3_6__14,linha3_6__13,linha3_6__12,linha3_6__11,linha3_6__10,
              linha3_6__9,linha3_6__8,linha3_6__7,linha3_6__6,linha3_6__5,
              linha3_6__4,linha3_6__3,linha3_6__2,linha3_6__1,linha3_6__0}), .a1 (
              {linha2_5__31,linha2_5__30,linha2_5__29,linha2_5__28,linha2_5__27,
              linha2_5__26,linha2_5__25,linha2_5__24,linha2_5__23,linha2_5__22,
              linha2_5__21,linha2_5__20,linha2_5__19,linha2_5__18,linha2_5__17,
              linha2_5__16,linha2_5__15,linha2_5__14,linha2_5__13,linha2_5__12,
              linha2_5__11,linha2_5__10,linha2_5__9,linha2_5__8,linha2_5__7,
              linha2_5__6,linha2_5__5,linha2_5__4,linha2_5__3,linha2_5__2,
              linha2_5__1,linha2_5__0}), .a0 ({linha3_5__31,linha3_5__30,
              linha3_5__29,linha3_5__28,linha3_5__27,linha3_5__26,linha3_5__25,
              linha3_5__24,linha3_5__23,linha3_5__22,linha3_5__21,linha3_5__20,
              linha3_5__19,linha3_5__18,linha3_5__17,linha3_5__16,linha3_5__15,
              linha3_5__14,linha3_5__13,linha3_5__12,linha3_5__11,linha3_5__10,
              linha3_5__9,linha3_5__8,linha3_5__7,linha3_5__6,linha3_5__5,
              linha3_5__4,linha3_5__3,linha3_5__2,linha3_5__1,linha3_5__0}), .s (
              row_5_rowi_bni1_l)) ;
    juntarComparadores_32 row_5_rowi_bni2_Comp (.g (\$dummy [19]), .l (
                          row_5_rowi_bni2_l), .a ({linha4_5__31,linha4_5__30,
                          linha4_5__29,linha4_5__28,linha4_5__27,linha4_5__26,
                          linha4_5__25,linha4_5__24,linha4_5__23,linha4_5__22,
                          linha4_5__21,linha4_5__20,linha4_5__19,linha4_5__18,
                          linha4_5__17,linha4_5__16,linha4_5__15,linha4_5__14,
                          linha4_5__13,linha4_5__12,linha4_5__11,linha4_5__10,
                          linha4_5__9,linha4_5__8,linha4_5__7,linha4_5__6,
                          linha4_5__5,linha4_5__4,linha4_5__3,linha4_5__2,
                          linha4_5__1,linha4_5__0}), .b ({linha5_5__31,
                          linha5_5__30,linha5_5__29,linha5_5__28,linha5_5__27,
                          linha5_5__26,linha5_5__25,linha5_5__24,linha5_5__23,
                          linha5_5__22,linha5_5__21,linha5_5__20,linha5_5__19,
                          linha5_5__18,linha5_5__17,linha5_5__16,linha5_5__15,
                          linha5_5__14,linha5_5__13,linha5_5__12,linha5_5__11,
                          linha5_5__10,linha5_5__9,linha5_5__8,linha5_5__7,
                          linha5_5__6,linha5_5__5,linha5_5__4,linha5_5__3,
                          linha5_5__2,linha5_5__1,linha5_5__0})) ;
    Mux2x1_32 row_5_rowi_bni2_muxMax (.r ({linha4_6__31,linha4_6__30,
              linha4_6__29,linha4_6__28,linha4_6__27,linha4_6__26,linha4_6__25,
              linha4_6__24,linha4_6__23,linha4_6__22,linha4_6__21,linha4_6__20,
              linha4_6__19,linha4_6__18,linha4_6__17,linha4_6__16,linha4_6__15,
              linha4_6__14,linha4_6__13,linha4_6__12,linha4_6__11,linha4_6__10,
              linha4_6__9,linha4_6__8,linha4_6__7,linha4_6__6,linha4_6__5,
              linha4_6__4,linha4_6__3,linha4_6__2,linha4_6__1,linha4_6__0}), .a1 (
              {linha5_5__31,linha5_5__30,linha5_5__29,linha5_5__28,linha5_5__27,
              linha5_5__26,linha5_5__25,linha5_5__24,linha5_5__23,linha5_5__22,
              linha5_5__21,linha5_5__20,linha5_5__19,linha5_5__18,linha5_5__17,
              linha5_5__16,linha5_5__15,linha5_5__14,linha5_5__13,linha5_5__12,
              linha5_5__11,linha5_5__10,linha5_5__9,linha5_5__8,linha5_5__7,
              linha5_5__6,linha5_5__5,linha5_5__4,linha5_5__3,linha5_5__2,
              linha5_5__1,linha5_5__0}), .a0 ({linha4_5__31,linha4_5__30,
              linha4_5__29,linha4_5__28,linha4_5__27,linha4_5__26,linha4_5__25,
              linha4_5__24,linha4_5__23,linha4_5__22,linha4_5__21,linha4_5__20,
              linha4_5__19,linha4_5__18,linha4_5__17,linha4_5__16,linha4_5__15,
              linha4_5__14,linha4_5__13,linha4_5__12,linha4_5__11,linha4_5__10,
              linha4_5__9,linha4_5__8,linha4_5__7,linha4_5__6,linha4_5__5,
              linha4_5__4,linha4_5__3,linha4_5__2,linha4_5__1,linha4_5__0}), .s (
              row_5_rowi_bni2_l)) ;
    Mux2x1_32 row_5_rowi_bni2_muxMin (.r ({linha5_6__31,linha5_6__30,
              linha5_6__29,linha5_6__28,linha5_6__27,linha5_6__26,linha5_6__25,
              linha5_6__24,linha5_6__23,linha5_6__22,linha5_6__21,linha5_6__20,
              linha5_6__19,linha5_6__18,linha5_6__17,linha5_6__16,linha5_6__15,
              linha5_6__14,linha5_6__13,linha5_6__12,linha5_6__11,linha5_6__10,
              linha5_6__9,linha5_6__8,linha5_6__7,linha5_6__6,linha5_6__5,
              linha5_6__4,linha5_6__3,linha5_6__2,linha5_6__1,linha5_6__0}), .a1 (
              {linha4_5__31,linha4_5__30,linha4_5__29,linha4_5__28,linha4_5__27,
              linha4_5__26,linha4_5__25,linha4_5__24,linha4_5__23,linha4_5__22,
              linha4_5__21,linha4_5__20,linha4_5__19,linha4_5__18,linha4_5__17,
              linha4_5__16,linha4_5__15,linha4_5__14,linha4_5__13,linha4_5__12,
              linha4_5__11,linha4_5__10,linha4_5__9,linha4_5__8,linha4_5__7,
              linha4_5__6,linha4_5__5,linha4_5__4,linha4_5__3,linha4_5__2,
              linha4_5__1,linha4_5__0}), .a0 ({linha5_5__31,linha5_5__30,
              linha5_5__29,linha5_5__28,linha5_5__27,linha5_5__26,linha5_5__25,
              linha5_5__24,linha5_5__23,linha5_5__22,linha5_5__21,linha5_5__20,
              linha5_5__19,linha5_5__18,linha5_5__17,linha5_5__16,linha5_5__15,
              linha5_5__14,linha5_5__13,linha5_5__12,linha5_5__11,linha5_5__10,
              linha5_5__9,linha5_5__8,linha5_5__7,linha5_5__6,linha5_5__5,
              linha5_5__4,linha5_5__3,linha5_5__2,linha5_5__1,linha5_5__0}), .s (
              row_5_rowi_bni2_l)) ;
    juntarComparadores_32 row_5_rowi_bni3_Comp (.g (\$dummy [20]), .l (
                          row_5_rowi_bni3_l), .a ({linha6_5__31,linha6_5__30,
                          linha6_5__29,linha6_5__28,linha6_5__27,linha6_5__26,
                          linha6_5__25,linha6_5__24,linha6_5__23,linha6_5__22,
                          linha6_5__21,linha6_5__20,linha6_5__19,linha6_5__18,
                          linha6_5__17,linha6_5__16,linha6_5__15,linha6_5__14,
                          linha6_5__13,linha6_5__12,linha6_5__11,linha6_5__10,
                          linha6_5__9,linha6_5__8,linha6_5__7,linha6_5__6,
                          linha6_5__5,linha6_5__4,linha6_5__3,linha6_5__2,
                          linha6_5__1,linha6_5__0}), .b ({linha7_5__31,
                          linha7_5__30,linha7_5__29,linha7_5__28,linha7_5__27,
                          linha7_5__26,linha7_5__25,linha7_5__24,linha7_5__23,
                          linha7_5__22,linha7_5__21,linha7_5__20,linha7_5__19,
                          linha7_5__18,linha7_5__17,linha7_5__16,linha7_5__15,
                          linha7_5__14,linha7_5__13,linha7_5__12,linha7_5__11,
                          linha7_5__10,linha7_5__9,linha7_5__8,linha7_5__7,
                          linha7_5__6,linha7_5__5,linha7_5__4,linha7_5__3,
                          linha7_5__2,linha7_5__1,linha7_5__0})) ;
    Mux2x1_32 row_5_rowi_bni3_muxMax (.r ({linha6_6__31,linha6_6__30,
              linha6_6__29,linha6_6__28,linha6_6__27,linha6_6__26,linha6_6__25,
              linha6_6__24,linha6_6__23,linha6_6__22,linha6_6__21,linha6_6__20,
              linha6_6__19,linha6_6__18,linha6_6__17,linha6_6__16,linha6_6__15,
              linha6_6__14,linha6_6__13,linha6_6__12,linha6_6__11,linha6_6__10,
              linha6_6__9,linha6_6__8,linha6_6__7,linha6_6__6,linha6_6__5,
              linha6_6__4,linha6_6__3,linha6_6__2,linha6_6__1,linha6_6__0}), .a1 (
              {linha7_5__31,linha7_5__30,linha7_5__29,linha7_5__28,linha7_5__27,
              linha7_5__26,linha7_5__25,linha7_5__24,linha7_5__23,linha7_5__22,
              linha7_5__21,linha7_5__20,linha7_5__19,linha7_5__18,linha7_5__17,
              linha7_5__16,linha7_5__15,linha7_5__14,linha7_5__13,linha7_5__12,
              linha7_5__11,linha7_5__10,linha7_5__9,linha7_5__8,linha7_5__7,
              linha7_5__6,linha7_5__5,linha7_5__4,linha7_5__3,linha7_5__2,
              linha7_5__1,linha7_5__0}), .a0 ({linha6_5__31,linha6_5__30,
              linha6_5__29,linha6_5__28,linha6_5__27,linha6_5__26,linha6_5__25,
              linha6_5__24,linha6_5__23,linha6_5__22,linha6_5__21,linha6_5__20,
              linha6_5__19,linha6_5__18,linha6_5__17,linha6_5__16,linha6_5__15,
              linha6_5__14,linha6_5__13,linha6_5__12,linha6_5__11,linha6_5__10,
              linha6_5__9,linha6_5__8,linha6_5__7,linha6_5__6,linha6_5__5,
              linha6_5__4,linha6_5__3,linha6_5__2,linha6_5__1,linha6_5__0}), .s (
              row_5_rowi_bni3_l)) ;
    Mux2x1_32 row_5_rowi_bni3_muxMin (.r ({linha7_6__31,linha7_6__30,
              linha7_6__29,linha7_6__28,linha7_6__27,linha7_6__26,linha7_6__25,
              linha7_6__24,linha7_6__23,linha7_6__22,linha7_6__21,linha7_6__20,
              linha7_6__19,linha7_6__18,linha7_6__17,linha7_6__16,linha7_6__15,
              linha7_6__14,linha7_6__13,linha7_6__12,linha7_6__11,linha7_6__10,
              linha7_6__9,linha7_6__8,linha7_6__7,linha7_6__6,linha7_6__5,
              linha7_6__4,linha7_6__3,linha7_6__2,linha7_6__1,linha7_6__0}), .a1 (
              {linha6_5__31,linha6_5__30,linha6_5__29,linha6_5__28,linha6_5__27,
              linha6_5__26,linha6_5__25,linha6_5__24,linha6_5__23,linha6_5__22,
              linha6_5__21,linha6_5__20,linha6_5__19,linha6_5__18,linha6_5__17,
              linha6_5__16,linha6_5__15,linha6_5__14,linha6_5__13,linha6_5__12,
              linha6_5__11,linha6_5__10,linha6_5__9,linha6_5__8,linha6_5__7,
              linha6_5__6,linha6_5__5,linha6_5__4,linha6_5__3,linha6_5__2,
              linha6_5__1,linha6_5__0}), .a0 ({linha7_5__31,linha7_5__30,
              linha7_5__29,linha7_5__28,linha7_5__27,linha7_5__26,linha7_5__25,
              linha7_5__24,linha7_5__23,linha7_5__22,linha7_5__21,linha7_5__20,
              linha7_5__19,linha7_5__18,linha7_5__17,linha7_5__16,linha7_5__15,
              linha7_5__14,linha7_5__13,linha7_5__12,linha7_5__11,linha7_5__10,
              linha7_5__9,linha7_5__8,linha7_5__7,linha7_5__6,linha7_5__5,
              linha7_5__4,linha7_5__3,linha7_5__2,linha7_5__1,linha7_5__0}), .s (
              row_5_rowi_bni3_l)) ;
    juntarComparadores_32 row_6_rowp_bni1_Comp (.g (\$dummy [21]), .l (
                          row_6_rowp_bni1_l), .a ({linha1_3__31,linha1_3__30,
                          linha1_3__29,linha1_3__28,linha1_3__27,linha1_3__26,
                          linha1_3__25,linha1_3__24,linha1_3__23,linha1_3__22,
                          linha1_3__21,linha1_3__20,linha1_3__19,linha1_3__18,
                          linha1_3__17,linha1_3__16,linha1_3__15,linha1_3__14,
                          linha1_3__13,linha1_3__12,linha1_3__11,linha1_3__10,
                          linha1_3__9,linha1_3__8,linha1_3__7,linha1_3__6,
                          linha1_3__5,linha1_3__4,linha1_3__3,linha1_3__2,
                          linha1_3__1,linha1_3__0}), .b ({linha2_6__31,
                          linha2_6__30,linha2_6__29,linha2_6__28,linha2_6__27,
                          linha2_6__26,linha2_6__25,linha2_6__24,linha2_6__23,
                          linha2_6__22,linha2_6__21,linha2_6__20,linha2_6__19,
                          linha2_6__18,linha2_6__17,linha2_6__16,linha2_6__15,
                          linha2_6__14,linha2_6__13,linha2_6__12,linha2_6__11,
                          linha2_6__10,linha2_6__9,linha2_6__8,linha2_6__7,
                          linha2_6__6,linha2_6__5,linha2_6__4,linha2_6__3,
                          linha2_6__2,linha2_6__1,linha2_6__0})) ;
    Mux2x1_32 row_6_rowp_bni1_muxMax (.r ({y1[31],y1[30],y1[29],y1[28],y1[27],
              y1[26],y1[25],y1[24],y1[23],y1[22],y1[21],y1[20],y1[19],y1[18],
              y1[17],y1[16],y1[15],y1[14],y1[13],y1[12],y1[11],y1[10],y1[9],
              y1[8],y1[7],y1[6],y1[5],y1[4],y1[3],y1[2],y1[1],y1[0]}), .a1 ({
              linha2_6__31,linha2_6__30,linha2_6__29,linha2_6__28,linha2_6__27,
              linha2_6__26,linha2_6__25,linha2_6__24,linha2_6__23,linha2_6__22,
              linha2_6__21,linha2_6__20,linha2_6__19,linha2_6__18,linha2_6__17,
              linha2_6__16,linha2_6__15,linha2_6__14,linha2_6__13,linha2_6__12,
              linha2_6__11,linha2_6__10,linha2_6__9,linha2_6__8,linha2_6__7,
              linha2_6__6,linha2_6__5,linha2_6__4,linha2_6__3,linha2_6__2,
              linha2_6__1,linha2_6__0}), .a0 ({linha1_3__31,linha1_3__30,
              linha1_3__29,linha1_3__28,linha1_3__27,linha1_3__26,linha1_3__25,
              linha1_3__24,linha1_3__23,linha1_3__22,linha1_3__21,linha1_3__20,
              linha1_3__19,linha1_3__18,linha1_3__17,linha1_3__16,linha1_3__15,
              linha1_3__14,linha1_3__13,linha1_3__12,linha1_3__11,linha1_3__10,
              linha1_3__9,linha1_3__8,linha1_3__7,linha1_3__6,linha1_3__5,
              linha1_3__4,linha1_3__3,linha1_3__2,linha1_3__1,linha1_3__0}), .s (
              row_6_rowp_bni1_l)) ;
    Mux2x1_32 row_6_rowp_bni1_muxMin (.r ({linha2_7__31,linha2_7__30,
              linha2_7__29,linha2_7__28,linha2_7__27,linha2_7__26,linha2_7__25,
              linha2_7__24,linha2_7__23,linha2_7__22,linha2_7__21,linha2_7__20,
              linha2_7__19,linha2_7__18,linha2_7__17,linha2_7__16,linha2_7__15,
              linha2_7__14,linha2_7__13,linha2_7__12,linha2_7__11,linha2_7__10,
              linha2_7__9,linha2_7__8,linha2_7__7,linha2_7__6,linha2_7__5,
              linha2_7__4,linha2_7__3,linha2_7__2,linha2_7__1,linha2_7__0}), .a1 (
              {linha1_3__31,linha1_3__30,linha1_3__29,linha1_3__28,linha1_3__27,
              linha1_3__26,linha1_3__25,linha1_3__24,linha1_3__23,linha1_3__22,
              linha1_3__21,linha1_3__20,linha1_3__19,linha1_3__18,linha1_3__17,
              linha1_3__16,linha1_3__15,linha1_3__14,linha1_3__13,linha1_3__12,
              linha1_3__11,linha1_3__10,linha1_3__9,linha1_3__8,linha1_3__7,
              linha1_3__6,linha1_3__5,linha1_3__4,linha1_3__3,linha1_3__2,
              linha1_3__1,linha1_3__0}), .a0 ({linha2_6__31,linha2_6__30,
              linha2_6__29,linha2_6__28,linha2_6__27,linha2_6__26,linha2_6__25,
              linha2_6__24,linha2_6__23,linha2_6__22,linha2_6__21,linha2_6__20,
              linha2_6__19,linha2_6__18,linha2_6__17,linha2_6__16,linha2_6__15,
              linha2_6__14,linha2_6__13,linha2_6__12,linha2_6__11,linha2_6__10,
              linha2_6__9,linha2_6__8,linha2_6__7,linha2_6__6,linha2_6__5,
              linha2_6__4,linha2_6__3,linha2_6__2,linha2_6__1,linha2_6__0}), .s (
              row_6_rowp_bni1_l)) ;
    juntarComparadores_32 row_6_rowp_bni2_Comp (.g (\$dummy [22]), .l (
                          row_6_rowp_bni2_l), .a ({linha3_6__31,linha3_6__30,
                          linha3_6__29,linha3_6__28,linha3_6__27,linha3_6__26,
                          linha3_6__25,linha3_6__24,linha3_6__23,linha3_6__22,
                          linha3_6__21,linha3_6__20,linha3_6__19,linha3_6__18,
                          linha3_6__17,linha3_6__16,linha3_6__15,linha3_6__14,
                          linha3_6__13,linha3_6__12,linha3_6__11,linha3_6__10,
                          linha3_6__9,linha3_6__8,linha3_6__7,linha3_6__6,
                          linha3_6__5,linha3_6__4,linha3_6__3,linha3_6__2,
                          linha3_6__1,linha3_6__0}), .b ({linha4_6__31,
                          linha4_6__30,linha4_6__29,linha4_6__28,linha4_6__27,
                          linha4_6__26,linha4_6__25,linha4_6__24,linha4_6__23,
                          linha4_6__22,linha4_6__21,linha4_6__20,linha4_6__19,
                          linha4_6__18,linha4_6__17,linha4_6__16,linha4_6__15,
                          linha4_6__14,linha4_6__13,linha4_6__12,linha4_6__11,
                          linha4_6__10,linha4_6__9,linha4_6__8,linha4_6__7,
                          linha4_6__6,linha4_6__5,linha4_6__4,linha4_6__3,
                          linha4_6__2,linha4_6__1,linha4_6__0})) ;
    Mux2x1_32 row_6_rowp_bni2_muxMax (.r ({linha3_7__31,linha3_7__30,
              linha3_7__29,linha3_7__28,linha3_7__27,linha3_7__26,linha3_7__25,
              linha3_7__24,linha3_7__23,linha3_7__22,linha3_7__21,linha3_7__20,
              linha3_7__19,linha3_7__18,linha3_7__17,linha3_7__16,linha3_7__15,
              linha3_7__14,linha3_7__13,linha3_7__12,linha3_7__11,linha3_7__10,
              linha3_7__9,linha3_7__8,linha3_7__7,linha3_7__6,linha3_7__5,
              linha3_7__4,linha3_7__3,linha3_7__2,linha3_7__1,linha3_7__0}), .a1 (
              {linha4_6__31,linha4_6__30,linha4_6__29,linha4_6__28,linha4_6__27,
              linha4_6__26,linha4_6__25,linha4_6__24,linha4_6__23,linha4_6__22,
              linha4_6__21,linha4_6__20,linha4_6__19,linha4_6__18,linha4_6__17,
              linha4_6__16,linha4_6__15,linha4_6__14,linha4_6__13,linha4_6__12,
              linha4_6__11,linha4_6__10,linha4_6__9,linha4_6__8,linha4_6__7,
              linha4_6__6,linha4_6__5,linha4_6__4,linha4_6__3,linha4_6__2,
              linha4_6__1,linha4_6__0}), .a0 ({linha3_6__31,linha3_6__30,
              linha3_6__29,linha3_6__28,linha3_6__27,linha3_6__26,linha3_6__25,
              linha3_6__24,linha3_6__23,linha3_6__22,linha3_6__21,linha3_6__20,
              linha3_6__19,linha3_6__18,linha3_6__17,linha3_6__16,linha3_6__15,
              linha3_6__14,linha3_6__13,linha3_6__12,linha3_6__11,linha3_6__10,
              linha3_6__9,linha3_6__8,linha3_6__7,linha3_6__6,linha3_6__5,
              linha3_6__4,linha3_6__3,linha3_6__2,linha3_6__1,linha3_6__0}), .s (
              row_6_rowp_bni2_l)) ;
    Mux2x1_32 row_6_rowp_bni2_muxMin (.r ({linha4_7__31,linha4_7__30,
              linha4_7__29,linha4_7__28,linha4_7__27,linha4_7__26,linha4_7__25,
              linha4_7__24,linha4_7__23,linha4_7__22,linha4_7__21,linha4_7__20,
              linha4_7__19,linha4_7__18,linha4_7__17,linha4_7__16,linha4_7__15,
              linha4_7__14,linha4_7__13,linha4_7__12,linha4_7__11,linha4_7__10,
              linha4_7__9,linha4_7__8,linha4_7__7,linha4_7__6,linha4_7__5,
              linha4_7__4,linha4_7__3,linha4_7__2,linha4_7__1,linha4_7__0}), .a1 (
              {linha3_6__31,linha3_6__30,linha3_6__29,linha3_6__28,linha3_6__27,
              linha3_6__26,linha3_6__25,linha3_6__24,linha3_6__23,linha3_6__22,
              linha3_6__21,linha3_6__20,linha3_6__19,linha3_6__18,linha3_6__17,
              linha3_6__16,linha3_6__15,linha3_6__14,linha3_6__13,linha3_6__12,
              linha3_6__11,linha3_6__10,linha3_6__9,linha3_6__8,linha3_6__7,
              linha3_6__6,linha3_6__5,linha3_6__4,linha3_6__3,linha3_6__2,
              linha3_6__1,linha3_6__0}), .a0 ({linha4_6__31,linha4_6__30,
              linha4_6__29,linha4_6__28,linha4_6__27,linha4_6__26,linha4_6__25,
              linha4_6__24,linha4_6__23,linha4_6__22,linha4_6__21,linha4_6__20,
              linha4_6__19,linha4_6__18,linha4_6__17,linha4_6__16,linha4_6__15,
              linha4_6__14,linha4_6__13,linha4_6__12,linha4_6__11,linha4_6__10,
              linha4_6__9,linha4_6__8,linha4_6__7,linha4_6__6,linha4_6__5,
              linha4_6__4,linha4_6__3,linha4_6__2,linha4_6__1,linha4_6__0}), .s (
              row_6_rowp_bni2_l)) ;
    juntarComparadores_32 row_6_rowp_bni3_Comp (.g (\$dummy [23]), .l (
                          row_6_rowp_bni3_l), .a ({linha5_6__31,linha5_6__30,
                          linha5_6__29,linha5_6__28,linha5_6__27,linha5_6__26,
                          linha5_6__25,linha5_6__24,linha5_6__23,linha5_6__22,
                          linha5_6__21,linha5_6__20,linha5_6__19,linha5_6__18,
                          linha5_6__17,linha5_6__16,linha5_6__15,linha5_6__14,
                          linha5_6__13,linha5_6__12,linha5_6__11,linha5_6__10,
                          linha5_6__9,linha5_6__8,linha5_6__7,linha5_6__6,
                          linha5_6__5,linha5_6__4,linha5_6__3,linha5_6__2,
                          linha5_6__1,linha5_6__0}), .b ({linha6_6__31,
                          linha6_6__30,linha6_6__29,linha6_6__28,linha6_6__27,
                          linha6_6__26,linha6_6__25,linha6_6__24,linha6_6__23,
                          linha6_6__22,linha6_6__21,linha6_6__20,linha6_6__19,
                          linha6_6__18,linha6_6__17,linha6_6__16,linha6_6__15,
                          linha6_6__14,linha6_6__13,linha6_6__12,linha6_6__11,
                          linha6_6__10,linha6_6__9,linha6_6__8,linha6_6__7,
                          linha6_6__6,linha6_6__5,linha6_6__4,linha6_6__3,
                          linha6_6__2,linha6_6__1,linha6_6__0})) ;
    Mux2x1_32 row_6_rowp_bni3_muxMax (.r ({linha5_7__31,linha5_7__30,
              linha5_7__29,linha5_7__28,linha5_7__27,linha5_7__26,linha5_7__25,
              linha5_7__24,linha5_7__23,linha5_7__22,linha5_7__21,linha5_7__20,
              linha5_7__19,linha5_7__18,linha5_7__17,linha5_7__16,linha5_7__15,
              linha5_7__14,linha5_7__13,linha5_7__12,linha5_7__11,linha5_7__10,
              linha5_7__9,linha5_7__8,linha5_7__7,linha5_7__6,linha5_7__5,
              linha5_7__4,linha5_7__3,linha5_7__2,linha5_7__1,linha5_7__0}), .a1 (
              {linha6_6__31,linha6_6__30,linha6_6__29,linha6_6__28,linha6_6__27,
              linha6_6__26,linha6_6__25,linha6_6__24,linha6_6__23,linha6_6__22,
              linha6_6__21,linha6_6__20,linha6_6__19,linha6_6__18,linha6_6__17,
              linha6_6__16,linha6_6__15,linha6_6__14,linha6_6__13,linha6_6__12,
              linha6_6__11,linha6_6__10,linha6_6__9,linha6_6__8,linha6_6__7,
              linha6_6__6,linha6_6__5,linha6_6__4,linha6_6__3,linha6_6__2,
              linha6_6__1,linha6_6__0}), .a0 ({linha5_6__31,linha5_6__30,
              linha5_6__29,linha5_6__28,linha5_6__27,linha5_6__26,linha5_6__25,
              linha5_6__24,linha5_6__23,linha5_6__22,linha5_6__21,linha5_6__20,
              linha5_6__19,linha5_6__18,linha5_6__17,linha5_6__16,linha5_6__15,
              linha5_6__14,linha5_6__13,linha5_6__12,linha5_6__11,linha5_6__10,
              linha5_6__9,linha5_6__8,linha5_6__7,linha5_6__6,linha5_6__5,
              linha5_6__4,linha5_6__3,linha5_6__2,linha5_6__1,linha5_6__0}), .s (
              row_6_rowp_bni3_l)) ;
    Mux2x1_32 row_6_rowp_bni3_muxMin (.r ({linha6_7__31,linha6_7__30,
              linha6_7__29,linha6_7__28,linha6_7__27,linha6_7__26,linha6_7__25,
              linha6_7__24,linha6_7__23,linha6_7__22,linha6_7__21,linha6_7__20,
              linha6_7__19,linha6_7__18,linha6_7__17,linha6_7__16,linha6_7__15,
              linha6_7__14,linha6_7__13,linha6_7__12,linha6_7__11,linha6_7__10,
              linha6_7__9,linha6_7__8,linha6_7__7,linha6_7__6,linha6_7__5,
              linha6_7__4,linha6_7__3,linha6_7__2,linha6_7__1,linha6_7__0}), .a1 (
              {linha5_6__31,linha5_6__30,linha5_6__29,linha5_6__28,linha5_6__27,
              linha5_6__26,linha5_6__25,linha5_6__24,linha5_6__23,linha5_6__22,
              linha5_6__21,linha5_6__20,linha5_6__19,linha5_6__18,linha5_6__17,
              linha5_6__16,linha5_6__15,linha5_6__14,linha5_6__13,linha5_6__12,
              linha5_6__11,linha5_6__10,linha5_6__9,linha5_6__8,linha5_6__7,
              linha5_6__6,linha5_6__5,linha5_6__4,linha5_6__3,linha5_6__2,
              linha5_6__1,linha5_6__0}), .a0 ({linha6_6__31,linha6_6__30,
              linha6_6__29,linha6_6__28,linha6_6__27,linha6_6__26,linha6_6__25,
              linha6_6__24,linha6_6__23,linha6_6__22,linha6_6__21,linha6_6__20,
              linha6_6__19,linha6_6__18,linha6_6__17,linha6_6__16,linha6_6__15,
              linha6_6__14,linha6_6__13,linha6_6__12,linha6_6__11,linha6_6__10,
              linha6_6__9,linha6_6__8,linha6_6__7,linha6_6__6,linha6_6__5,
              linha6_6__4,linha6_6__3,linha6_6__2,linha6_6__1,linha6_6__0}), .s (
              row_6_rowp_bni3_l)) ;
    juntarComparadores_32 row_6_rowp_bni4_Comp (.g (\$dummy [24]), .l (
                          row_6_rowp_bni4_l), .a ({linha7_6__31,linha7_6__30,
                          linha7_6__29,linha7_6__28,linha7_6__27,linha7_6__26,
                          linha7_6__25,linha7_6__24,linha7_6__23,linha7_6__22,
                          linha7_6__21,linha7_6__20,linha7_6__19,linha7_6__18,
                          linha7_6__17,linha7_6__16,linha7_6__15,linha7_6__14,
                          linha7_6__13,linha7_6__12,linha7_6__11,linha7_6__10,
                          linha7_6__9,linha7_6__8,linha7_6__7,linha7_6__6,
                          linha7_6__5,linha7_6__4,linha7_6__3,linha7_6__2,
                          linha7_6__1,linha7_6__0}), .b ({linha8_3__31,
                          linha8_3__30,linha8_3__29,linha8_3__28,linha8_3__27,
                          linha8_3__26,linha8_3__25,linha8_3__24,linha8_3__23,
                          linha8_3__22,linha8_3__21,linha8_3__20,linha8_3__19,
                          linha8_3__18,linha8_3__17,linha8_3__16,linha8_3__15,
                          linha8_3__14,linha8_3__13,linha8_3__12,linha8_3__11,
                          linha8_3__10,linha8_3__9,linha8_3__8,linha8_3__7,
                          linha8_3__6,linha8_3__5,linha8_3__4,linha8_3__3,
                          linha8_3__2,linha8_3__1,linha8_3__0})) ;
    Mux2x1_32 row_6_rowp_bni4_muxMax (.r ({linha7_7__31,linha7_7__30,
              linha7_7__29,linha7_7__28,linha7_7__27,linha7_7__26,linha7_7__25,
              linha7_7__24,linha7_7__23,linha7_7__22,linha7_7__21,linha7_7__20,
              linha7_7__19,linha7_7__18,linha7_7__17,linha7_7__16,linha7_7__15,
              linha7_7__14,linha7_7__13,linha7_7__12,linha7_7__11,linha7_7__10,
              linha7_7__9,linha7_7__8,linha7_7__7,linha7_7__6,linha7_7__5,
              linha7_7__4,linha7_7__3,linha7_7__2,linha7_7__1,linha7_7__0}), .a1 (
              {linha8_3__31,linha8_3__30,linha8_3__29,linha8_3__28,linha8_3__27,
              linha8_3__26,linha8_3__25,linha8_3__24,linha8_3__23,linha8_3__22,
              linha8_3__21,linha8_3__20,linha8_3__19,linha8_3__18,linha8_3__17,
              linha8_3__16,linha8_3__15,linha8_3__14,linha8_3__13,linha8_3__12,
              linha8_3__11,linha8_3__10,linha8_3__9,linha8_3__8,linha8_3__7,
              linha8_3__6,linha8_3__5,linha8_3__4,linha8_3__3,linha8_3__2,
              linha8_3__1,linha8_3__0}), .a0 ({linha7_6__31,linha7_6__30,
              linha7_6__29,linha7_6__28,linha7_6__27,linha7_6__26,linha7_6__25,
              linha7_6__24,linha7_6__23,linha7_6__22,linha7_6__21,linha7_6__20,
              linha7_6__19,linha7_6__18,linha7_6__17,linha7_6__16,linha7_6__15,
              linha7_6__14,linha7_6__13,linha7_6__12,linha7_6__11,linha7_6__10,
              linha7_6__9,linha7_6__8,linha7_6__7,linha7_6__6,linha7_6__5,
              linha7_6__4,linha7_6__3,linha7_6__2,linha7_6__1,linha7_6__0}), .s (
              row_6_rowp_bni4_l)) ;
    Mux2x1_32 row_6_rowp_bni4_muxMin (.r ({y8[31],y8[30],y8[29],y8[28],y8[27],
              y8[26],y8[25],y8[24],y8[23],y8[22],y8[21],y8[20],y8[19],y8[18],
              y8[17],y8[16],y8[15],y8[14],y8[13],y8[12],y8[11],y8[10],y8[9],
              y8[8],y8[7],y8[6],y8[5],y8[4],y8[3],y8[2],y8[1],y8[0]}), .a1 ({
              linha7_6__31,linha7_6__30,linha7_6__29,linha7_6__28,linha7_6__27,
              linha7_6__26,linha7_6__25,linha7_6__24,linha7_6__23,linha7_6__22,
              linha7_6__21,linha7_6__20,linha7_6__19,linha7_6__18,linha7_6__17,
              linha7_6__16,linha7_6__15,linha7_6__14,linha7_6__13,linha7_6__12,
              linha7_6__11,linha7_6__10,linha7_6__9,linha7_6__8,linha7_6__7,
              linha7_6__6,linha7_6__5,linha7_6__4,linha7_6__3,linha7_6__2,
              linha7_6__1,linha7_6__0}), .a0 ({linha8_3__31,linha8_3__30,
              linha8_3__29,linha8_3__28,linha8_3__27,linha8_3__26,linha8_3__25,
              linha8_3__24,linha8_3__23,linha8_3__22,linha8_3__21,linha8_3__20,
              linha8_3__19,linha8_3__18,linha8_3__17,linha8_3__16,linha8_3__15,
              linha8_3__14,linha8_3__13,linha8_3__12,linha8_3__11,linha8_3__10,
              linha8_3__9,linha8_3__8,linha8_3__7,linha8_3__6,linha8_3__5,
              linha8_3__4,linha8_3__3,linha8_3__2,linha8_3__1,linha8_3__0}), .s (
              row_6_rowp_bni4_l)) ;
    juntarComparadores_32 row_7_rowi_bni1_Comp (.g (\$dummy [25]), .l (
                          row_7_rowi_bni1_l), .a ({linha2_7__31,linha2_7__30,
                          linha2_7__29,linha2_7__28,linha2_7__27,linha2_7__26,
                          linha2_7__25,linha2_7__24,linha2_7__23,linha2_7__22,
                          linha2_7__21,linha2_7__20,linha2_7__19,linha2_7__18,
                          linha2_7__17,linha2_7__16,linha2_7__15,linha2_7__14,
                          linha2_7__13,linha2_7__12,linha2_7__11,linha2_7__10,
                          linha2_7__9,linha2_7__8,linha2_7__7,linha2_7__6,
                          linha2_7__5,linha2_7__4,linha2_7__3,linha2_7__2,
                          linha2_7__1,linha2_7__0}), .b ({linha3_7__31,
                          linha3_7__30,linha3_7__29,linha3_7__28,linha3_7__27,
                          linha3_7__26,linha3_7__25,linha3_7__24,linha3_7__23,
                          linha3_7__22,linha3_7__21,linha3_7__20,linha3_7__19,
                          linha3_7__18,linha3_7__17,linha3_7__16,linha3_7__15,
                          linha3_7__14,linha3_7__13,linha3_7__12,linha3_7__11,
                          linha3_7__10,linha3_7__9,linha3_7__8,linha3_7__7,
                          linha3_7__6,linha3_7__5,linha3_7__4,linha3_7__3,
                          linha3_7__2,linha3_7__1,linha3_7__0})) ;
    Mux2x1_32 row_7_rowi_bni1_muxMax (.r ({y2[31],y2[30],y2[29],y2[28],y2[27],
              y2[26],y2[25],y2[24],y2[23],y2[22],y2[21],y2[20],y2[19],y2[18],
              y2[17],y2[16],y2[15],y2[14],y2[13],y2[12],y2[11],y2[10],y2[9],
              y2[8],y2[7],y2[6],y2[5],y2[4],y2[3],y2[2],y2[1],y2[0]}), .a1 ({
              linha3_7__31,linha3_7__30,linha3_7__29,linha3_7__28,linha3_7__27,
              linha3_7__26,linha3_7__25,linha3_7__24,linha3_7__23,linha3_7__22,
              linha3_7__21,linha3_7__20,linha3_7__19,linha3_7__18,linha3_7__17,
              linha3_7__16,linha3_7__15,linha3_7__14,linha3_7__13,linha3_7__12,
              linha3_7__11,linha3_7__10,linha3_7__9,linha3_7__8,linha3_7__7,
              linha3_7__6,linha3_7__5,linha3_7__4,linha3_7__3,linha3_7__2,
              linha3_7__1,linha3_7__0}), .a0 ({linha2_7__31,linha2_7__30,
              linha2_7__29,linha2_7__28,linha2_7__27,linha2_7__26,linha2_7__25,
              linha2_7__24,linha2_7__23,linha2_7__22,linha2_7__21,linha2_7__20,
              linha2_7__19,linha2_7__18,linha2_7__17,linha2_7__16,linha2_7__15,
              linha2_7__14,linha2_7__13,linha2_7__12,linha2_7__11,linha2_7__10,
              linha2_7__9,linha2_7__8,linha2_7__7,linha2_7__6,linha2_7__5,
              linha2_7__4,linha2_7__3,linha2_7__2,linha2_7__1,linha2_7__0}), .s (
              row_7_rowi_bni1_l)) ;
    Mux2x1_32 row_7_rowi_bni1_muxMin (.r ({y3[31],y3[30],y3[29],y3[28],y3[27],
              y3[26],y3[25],y3[24],y3[23],y3[22],y3[21],y3[20],y3[19],y3[18],
              y3[17],y3[16],y3[15],y3[14],y3[13],y3[12],y3[11],y3[10],y3[9],
              y3[8],y3[7],y3[6],y3[5],y3[4],y3[3],y3[2],y3[1],y3[0]}), .a1 ({
              linha2_7__31,linha2_7__30,linha2_7__29,linha2_7__28,linha2_7__27,
              linha2_7__26,linha2_7__25,linha2_7__24,linha2_7__23,linha2_7__22,
              linha2_7__21,linha2_7__20,linha2_7__19,linha2_7__18,linha2_7__17,
              linha2_7__16,linha2_7__15,linha2_7__14,linha2_7__13,linha2_7__12,
              linha2_7__11,linha2_7__10,linha2_7__9,linha2_7__8,linha2_7__7,
              linha2_7__6,linha2_7__5,linha2_7__4,linha2_7__3,linha2_7__2,
              linha2_7__1,linha2_7__0}), .a0 ({linha3_7__31,linha3_7__30,
              linha3_7__29,linha3_7__28,linha3_7__27,linha3_7__26,linha3_7__25,
              linha3_7__24,linha3_7__23,linha3_7__22,linha3_7__21,linha3_7__20,
              linha3_7__19,linha3_7__18,linha3_7__17,linha3_7__16,linha3_7__15,
              linha3_7__14,linha3_7__13,linha3_7__12,linha3_7__11,linha3_7__10,
              linha3_7__9,linha3_7__8,linha3_7__7,linha3_7__6,linha3_7__5,
              linha3_7__4,linha3_7__3,linha3_7__2,linha3_7__1,linha3_7__0}), .s (
              row_7_rowi_bni1_l)) ;
    juntarComparadores_32 row_7_rowi_bni2_Comp (.g (\$dummy [26]), .l (
                          row_7_rowi_bni2_l), .a ({linha4_7__31,linha4_7__30,
                          linha4_7__29,linha4_7__28,linha4_7__27,linha4_7__26,
                          linha4_7__25,linha4_7__24,linha4_7__23,linha4_7__22,
                          linha4_7__21,linha4_7__20,linha4_7__19,linha4_7__18,
                          linha4_7__17,linha4_7__16,linha4_7__15,linha4_7__14,
                          linha4_7__13,linha4_7__12,linha4_7__11,linha4_7__10,
                          linha4_7__9,linha4_7__8,linha4_7__7,linha4_7__6,
                          linha4_7__5,linha4_7__4,linha4_7__3,linha4_7__2,
                          linha4_7__1,linha4_7__0}), .b ({linha5_7__31,
                          linha5_7__30,linha5_7__29,linha5_7__28,linha5_7__27,
                          linha5_7__26,linha5_7__25,linha5_7__24,linha5_7__23,
                          linha5_7__22,linha5_7__21,linha5_7__20,linha5_7__19,
                          linha5_7__18,linha5_7__17,linha5_7__16,linha5_7__15,
                          linha5_7__14,linha5_7__13,linha5_7__12,linha5_7__11,
                          linha5_7__10,linha5_7__9,linha5_7__8,linha5_7__7,
                          linha5_7__6,linha5_7__5,linha5_7__4,linha5_7__3,
                          linha5_7__2,linha5_7__1,linha5_7__0})) ;
    Mux2x1_32 row_7_rowi_bni2_muxMax (.r ({y4[31],y4[30],y4[29],y4[28],y4[27],
              y4[26],y4[25],y4[24],y4[23],y4[22],y4[21],y4[20],y4[19],y4[18],
              y4[17],y4[16],y4[15],y4[14],y4[13],y4[12],y4[11],y4[10],y4[9],
              y4[8],y4[7],y4[6],y4[5],y4[4],y4[3],y4[2],y4[1],y4[0]}), .a1 ({
              linha5_7__31,linha5_7__30,linha5_7__29,linha5_7__28,linha5_7__27,
              linha5_7__26,linha5_7__25,linha5_7__24,linha5_7__23,linha5_7__22,
              linha5_7__21,linha5_7__20,linha5_7__19,linha5_7__18,linha5_7__17,
              linha5_7__16,linha5_7__15,linha5_7__14,linha5_7__13,linha5_7__12,
              linha5_7__11,linha5_7__10,linha5_7__9,linha5_7__8,linha5_7__7,
              linha5_7__6,linha5_7__5,linha5_7__4,linha5_7__3,linha5_7__2,
              linha5_7__1,linha5_7__0}), .a0 ({linha4_7__31,linha4_7__30,
              linha4_7__29,linha4_7__28,linha4_7__27,linha4_7__26,linha4_7__25,
              linha4_7__24,linha4_7__23,linha4_7__22,linha4_7__21,linha4_7__20,
              linha4_7__19,linha4_7__18,linha4_7__17,linha4_7__16,linha4_7__15,
              linha4_7__14,linha4_7__13,linha4_7__12,linha4_7__11,linha4_7__10,
              linha4_7__9,linha4_7__8,linha4_7__7,linha4_7__6,linha4_7__5,
              linha4_7__4,linha4_7__3,linha4_7__2,linha4_7__1,linha4_7__0}), .s (
              row_7_rowi_bni2_l)) ;
    Mux2x1_32 row_7_rowi_bni2_muxMin (.r ({y5[31],y5[30],y5[29],y5[28],y5[27],
              y5[26],y5[25],y5[24],y5[23],y5[22],y5[21],y5[20],y5[19],y5[18],
              y5[17],y5[16],y5[15],y5[14],y5[13],y5[12],y5[11],y5[10],y5[9],
              y5[8],y5[7],y5[6],y5[5],y5[4],y5[3],y5[2],y5[1],y5[0]}), .a1 ({
              linha4_7__31,linha4_7__30,linha4_7__29,linha4_7__28,linha4_7__27,
              linha4_7__26,linha4_7__25,linha4_7__24,linha4_7__23,linha4_7__22,
              linha4_7__21,linha4_7__20,linha4_7__19,linha4_7__18,linha4_7__17,
              linha4_7__16,linha4_7__15,linha4_7__14,linha4_7__13,linha4_7__12,
              linha4_7__11,linha4_7__10,linha4_7__9,linha4_7__8,linha4_7__7,
              linha4_7__6,linha4_7__5,linha4_7__4,linha4_7__3,linha4_7__2,
              linha4_7__1,linha4_7__0}), .a0 ({linha5_7__31,linha5_7__30,
              linha5_7__29,linha5_7__28,linha5_7__27,linha5_7__26,linha5_7__25,
              linha5_7__24,linha5_7__23,linha5_7__22,linha5_7__21,linha5_7__20,
              linha5_7__19,linha5_7__18,linha5_7__17,linha5_7__16,linha5_7__15,
              linha5_7__14,linha5_7__13,linha5_7__12,linha5_7__11,linha5_7__10,
              linha5_7__9,linha5_7__8,linha5_7__7,linha5_7__6,linha5_7__5,
              linha5_7__4,linha5_7__3,linha5_7__2,linha5_7__1,linha5_7__0}), .s (
              row_7_rowi_bni2_l)) ;
    juntarComparadores_32 row_7_rowi_bni3_Comp (.g (\$dummy [27]), .l (
                          row_7_rowi_bni3_l), .a ({linha6_7__31,linha6_7__30,
                          linha6_7__29,linha6_7__28,linha6_7__27,linha6_7__26,
                          linha6_7__25,linha6_7__24,linha6_7__23,linha6_7__22,
                          linha6_7__21,linha6_7__20,linha6_7__19,linha6_7__18,
                          linha6_7__17,linha6_7__16,linha6_7__15,linha6_7__14,
                          linha6_7__13,linha6_7__12,linha6_7__11,linha6_7__10,
                          linha6_7__9,linha6_7__8,linha6_7__7,linha6_7__6,
                          linha6_7__5,linha6_7__4,linha6_7__3,linha6_7__2,
                          linha6_7__1,linha6_7__0}), .b ({linha7_7__31,
                          linha7_7__30,linha7_7__29,linha7_7__28,linha7_7__27,
                          linha7_7__26,linha7_7__25,linha7_7__24,linha7_7__23,
                          linha7_7__22,linha7_7__21,linha7_7__20,linha7_7__19,
                          linha7_7__18,linha7_7__17,linha7_7__16,linha7_7__15,
                          linha7_7__14,linha7_7__13,linha7_7__12,linha7_7__11,
                          linha7_7__10,linha7_7__9,linha7_7__8,linha7_7__7,
                          linha7_7__6,linha7_7__5,linha7_7__4,linha7_7__3,
                          linha7_7__2,linha7_7__1,linha7_7__0})) ;
    Mux2x1_32 row_7_rowi_bni3_muxMax (.r ({y6[31],y6[30],y6[29],y6[28],y6[27],
              y6[26],y6[25],y6[24],y6[23],y6[22],y6[21],y6[20],y6[19],y6[18],
              y6[17],y6[16],y6[15],y6[14],y6[13],y6[12],y6[11],y6[10],y6[9],
              y6[8],y6[7],y6[6],y6[5],y6[4],y6[3],y6[2],y6[1],y6[0]}), .a1 ({
              linha7_7__31,linha7_7__30,linha7_7__29,linha7_7__28,linha7_7__27,
              linha7_7__26,linha7_7__25,linha7_7__24,linha7_7__23,linha7_7__22,
              linha7_7__21,linha7_7__20,linha7_7__19,linha7_7__18,linha7_7__17,
              linha7_7__16,linha7_7__15,linha7_7__14,linha7_7__13,linha7_7__12,
              linha7_7__11,linha7_7__10,linha7_7__9,linha7_7__8,linha7_7__7,
              linha7_7__6,linha7_7__5,linha7_7__4,linha7_7__3,linha7_7__2,
              linha7_7__1,linha7_7__0}), .a0 ({linha6_7__31,linha6_7__30,
              linha6_7__29,linha6_7__28,linha6_7__27,linha6_7__26,linha6_7__25,
              linha6_7__24,linha6_7__23,linha6_7__22,linha6_7__21,linha6_7__20,
              linha6_7__19,linha6_7__18,linha6_7__17,linha6_7__16,linha6_7__15,
              linha6_7__14,linha6_7__13,linha6_7__12,linha6_7__11,linha6_7__10,
              linha6_7__9,linha6_7__8,linha6_7__7,linha6_7__6,linha6_7__5,
              linha6_7__4,linha6_7__3,linha6_7__2,linha6_7__1,linha6_7__0}), .s (
              row_7_rowi_bni3_l)) ;
    Mux2x1_32 row_7_rowi_bni3_muxMin (.r ({y7[31],y7[30],y7[29],y7[28],y7[27],
              y7[26],y7[25],y7[24],y7[23],y7[22],y7[21],y7[20],y7[19],y7[18],
              y7[17],y7[16],y7[15],y7[14],y7[13],y7[12],y7[11],y7[10],y7[9],
              y7[8],y7[7],y7[6],y7[5],y7[4],y7[3],y7[2],y7[1],y7[0]}), .a1 ({
              linha6_7__31,linha6_7__30,linha6_7__29,linha6_7__28,linha6_7__27,
              linha6_7__26,linha6_7__25,linha6_7__24,linha6_7__23,linha6_7__22,
              linha6_7__21,linha6_7__20,linha6_7__19,linha6_7__18,linha6_7__17,
              linha6_7__16,linha6_7__15,linha6_7__14,linha6_7__13,linha6_7__12,
              linha6_7__11,linha6_7__10,linha6_7__9,linha6_7__8,linha6_7__7,
              linha6_7__6,linha6_7__5,linha6_7__4,linha6_7__3,linha6_7__2,
              linha6_7__1,linha6_7__0}), .a0 ({linha7_7__31,linha7_7__30,
              linha7_7__29,linha7_7__28,linha7_7__27,linha7_7__26,linha7_7__25,
              linha7_7__24,linha7_7__23,linha7_7__22,linha7_7__21,linha7_7__20,
              linha7_7__19,linha7_7__18,linha7_7__17,linha7_7__16,linha7_7__15,
              linha7_7__14,linha7_7__13,linha7_7__12,linha7_7__11,linha7_7__10,
              linha7_7__9,linha7_7__8,linha7_7__7,linha7_7__6,linha7_7__5,
              linha7_7__4,linha7_7__3,linha7_7__2,linha7_7__1,linha7_7__0}), .s (
              row_7_rowi_bni3_l)) ;
    AN1T0 ix4094 (.X (nx4095), .A (row_0_rowp_bni1_l)) ;
endmodule


module AN1T0 ( X, A ) ;

    output X ;
    input A ;




    assign X = A ;
endmodule


module Mux2x1_32 ( r, a1, a0, s ) ;

    output [31:0]r ;
    input [31:0]a1 ;
    input [31:0]a0 ;
    input s ;

    wire nx351;



    MX2T0 ix7 (.X (r[0]), .A (a1[0]), .B (a0[0]), .S (nx351)) ;
    MX2T0 ix15 (.X (r[1]), .A (a1[1]), .B (a0[1]), .S (nx351)) ;
    MX2T0 ix23 (.X (r[2]), .A (a1[2]), .B (a0[2]), .S (nx351)) ;
    MX2T0 ix31 (.X (r[3]), .A (a1[3]), .B (a0[3]), .S (nx351)) ;
    MX2T0 ix39 (.X (r[4]), .A (a1[4]), .B (a0[4]), .S (nx351)) ;
    MX2T0 ix47 (.X (r[5]), .A (a1[5]), .B (a0[5]), .S (nx351)) ;
    MX2T0 ix55 (.X (r[6]), .A (a1[6]), .B (a0[6]), .S (nx351)) ;
    MX2T0 ix63 (.X (r[7]), .A (a1[7]), .B (a0[7]), .S (nx351)) ;
    MX2T0 ix71 (.X (r[8]), .A (a1[8]), .B (a0[8]), .S (nx351)) ;
    MX2T0 ix79 (.X (r[9]), .A (a1[9]), .B (a0[9]), .S (nx351)) ;
    MX2T0 ix87 (.X (r[10]), .A (a1[10]), .B (a0[10]), .S (nx351)) ;
    MX2T0 ix95 (.X (r[11]), .A (a1[11]), .B (a0[11]), .S (nx351)) ;
    MX2T0 ix103 (.X (r[12]), .A (a1[12]), .B (a0[12]), .S (nx351)) ;
    MX2T0 ix111 (.X (r[13]), .A (a1[13]), .B (a0[13]), .S (nx351)) ;
    MX2T0 ix119 (.X (r[14]), .A (a1[14]), .B (a0[14]), .S (nx351)) ;
    MX2T0 ix127 (.X (r[15]), .A (a1[15]), .B (a0[15]), .S (nx351)) ;
    MX2T0 ix135 (.X (r[16]), .A (a1[16]), .B (a0[16]), .S (nx351)) ;
    MX2T0 ix143 (.X (r[17]), .A (a1[17]), .B (a0[17]), .S (nx351)) ;
    MX2T0 ix151 (.X (r[18]), .A (a1[18]), .B (a0[18]), .S (nx351)) ;
    MX2T0 ix159 (.X (r[19]), .A (a1[19]), .B (a0[19]), .S (nx351)) ;
    MX2T0 ix167 (.X (r[20]), .A (a1[20]), .B (a0[20]), .S (nx351)) ;
    MX2T0 ix175 (.X (r[21]), .A (a1[21]), .B (a0[21]), .S (nx351)) ;
    MX2T0 ix183 (.X (r[22]), .A (a1[22]), .B (a0[22]), .S (nx351)) ;
    MX2T0 ix191 (.X (r[23]), .A (a1[23]), .B (a0[23]), .S (nx351)) ;
    MX2T0 ix199 (.X (r[24]), .A (a1[24]), .B (a0[24]), .S (nx351)) ;
    MX2T0 ix207 (.X (r[25]), .A (a1[25]), .B (a0[25]), .S (nx351)) ;
    MX2T0 ix215 (.X (r[26]), .A (a1[26]), .B (a0[26]), .S (nx351)) ;
    MX2T0 ix223 (.X (r[27]), .A (a1[27]), .B (a0[27]), .S (nx351)) ;
    MX2T0 ix231 (.X (r[28]), .A (a1[28]), .B (a0[28]), .S (nx351)) ;
    MX2T0 ix239 (.X (r[29]), .A (a1[29]), .B (a0[29]), .S (nx351)) ;
    MX2T0 ix247 (.X (r[30]), .A (a1[30]), .B (a0[30]), .S (nx351)) ;
    MX2T0 ix255 (.X (r[31]), .A (a1[31]), .B (a0[31]), .S (nx351)) ;
    AN1V1 ix350 (.X (nx351), .A (s)) ;
endmodule


module AN1V1 ( X, A ) ;

    output X ;
    input A ;




    assign X = A ;
endmodule


module MX2T0 ( X, A, B, S ) ;

    output X ;
    input A ;
    input B ;
    input S ;

    wire NOT_S, nx2, nx4;



    assign NOT_S = ~S ;
    and (nx2, B, NOT_S) ;
    and (nx4, A, S) ;
    or (X, nx2, nx4) ;
endmodule


module juntarComparadores_32 ( g, l, a, b ) ;

    output g ;
    output l ;
    input [31:0]a ;
    input [31:0]b ;

    wire nx28, nx48, nx58, nx88, nx98, nx128, nx138, nx168, nx178, nx208, nx218, 
         nx248, nx258, nx288, nx298, nx328, nx338, nx368, nx378, nx408, nx418, 
         nx448, nx458, nx488, nx498, nx528, nx538, nx568, nx578, nx598, nx608, 
         nx491, nx493, nx495, nx497, nx499, nx501, nx503, nx505, nx507, nx509, 
         nx511, nx513, nx515, nx517, nx519, nx521, nx523, nx525, nx527, nx529, 
         nx531, nx533, nx535, nx537, nx539, nx541, nx543, nx545, nx547, nx549, 
         nx551, nx553, nx555, nx557, nx559, nx561, nx563, nx565, nx567, nx569, 
         nx571, nx573, nx575, nx577, nx579, nx581, nx583, nx585, nx587, nx589, 
         nx591, nx593, nx595, nx597, nx599, nx601, nx603, nx605, nx607, nx609, 
         nx611, nx613, nx615, nx617, nx619, nx621, nx774, nx776;



    OAI3R1 ix619 (.X (l), .A1 (nx608), .A2 (a[0]), .A3 (nx619), .B (nx621)) ;
    OAI3R1 ix609 (.X (nx608), .A1 (nx578), .A2 (nx615), .A3 (b[1]), .B (nx617)
           ) ;
    OAI3R1 ix579 (.X (nx578), .A1 (nx568), .A2 (a[2]), .A3 (nx611), .B (nx613)
           ) ;
    OAI3R1 ix569 (.X (nx568), .A1 (nx538), .A2 (nx607), .A3 (b[3]), .B (nx609)
           ) ;
    OAI3R1 ix539 (.X (nx538), .A1 (nx528), .A2 (a[4]), .A3 (nx603), .B (nx605)
           ) ;
    OAI3R1 ix529 (.X (nx528), .A1 (nx498), .A2 (nx599), .A3 (b[5]), .B (nx601)
           ) ;
    OAI3R1 ix499 (.X (nx498), .A1 (nx488), .A2 (a[6]), .A3 (nx595), .B (nx597)
           ) ;
    OAI3R0 ix489 (.X (nx488), .A1 (nx458), .A2 (nx591), .A3 (b[7]), .B (nx593)
           ) ;
    OAI3R0 ix459 (.X (nx458), .A1 (nx448), .A2 (a[8]), .A3 (nx587), .B (nx589)
           ) ;
    OAI3R0 ix449 (.X (nx448), .A1 (nx418), .A2 (nx583), .A3 (b[9]), .B (nx585)
           ) ;
    OAI3R0 ix419 (.X (nx418), .A1 (nx408), .A2 (a[10]), .A3 (nx579), .B (nx581)
           ) ;
    OAI3R0 ix409 (.X (nx408), .A1 (nx378), .A2 (nx575), .A3 (b[11]), .B (nx577)
           ) ;
    OAI3R0 ix379 (.X (nx378), .A1 (nx368), .A2 (a[12]), .A3 (nx571), .B (nx573)
           ) ;
    OAI3R0 ix369 (.X (nx368), .A1 (nx338), .A2 (nx567), .A3 (b[13]), .B (nx569)
           ) ;
    OAI3R0 ix339 (.X (nx338), .A1 (nx328), .A2 (a[14]), .A3 (nx563), .B (nx565)
           ) ;
    OAI3R0 ix329 (.X (nx328), .A1 (nx298), .A2 (nx559), .A3 (b[15]), .B (nx561)
           ) ;
    OAI3R0 ix299 (.X (nx298), .A1 (nx288), .A2 (a[16]), .A3 (nx555), .B (nx557)
           ) ;
    OAI3R0 ix289 (.X (nx288), .A1 (nx258), .A2 (nx551), .A3 (b[17]), .B (nx553)
           ) ;
    OAI3R0 ix259 (.X (nx258), .A1 (nx248), .A2 (a[18]), .A3 (nx547), .B (nx549)
           ) ;
    OAI3R0 ix249 (.X (nx248), .A1 (nx218), .A2 (nx543), .A3 (b[19]), .B (nx545)
           ) ;
    OAI3R0 ix219 (.X (nx218), .A1 (nx208), .A2 (a[20]), .A3 (nx539), .B (nx541)
           ) ;
    OAI3R0 ix209 (.X (nx208), .A1 (nx178), .A2 (nx535), .A3 (b[21]), .B (nx537)
           ) ;
    OAI3R0 ix179 (.X (nx178), .A1 (nx168), .A2 (a[22]), .A3 (nx531), .B (nx533)
           ) ;
    OAI3R0 ix169 (.X (nx168), .A1 (nx138), .A2 (nx527), .A3 (b[23]), .B (nx529)
           ) ;
    OAI3R0 ix139 (.X (nx138), .A1 (nx128), .A2 (a[24]), .A3 (nx523), .B (nx525)
           ) ;
    OAI3R0 ix129 (.X (nx128), .A1 (nx98), .A2 (nx519), .A3 (b[25]), .B (nx521)
           ) ;
    OAI3R0 ix99 (.X (nx98), .A1 (nx88), .A2 (a[26]), .A3 (nx515), .B (nx517)) ;
    OAI3R0 ix89 (.X (nx88), .A1 (nx58), .A2 (nx511), .A3 (b[27]), .B (nx513)) ;
    OAI3R0 ix59 (.X (nx58), .A1 (nx48), .A2 (a[28]), .A3 (nx507), .B (nx509)) ;
    OAI3R0 ix49 (.X (nx48), .A1 (nx28), .A2 (nx499), .A3 (b[29]), .B (nx501)) ;
    OAI1A0 ix29 (.X (nx28), .A1 (a[31]), .A2 (nx491), .B (nx493)) ;
    IV1N0 ix492 (.X (nx491), .A (b[31])) ;
    OAI3N0 ix494 (.X (nx493), .A1 (nx495), .A2 (b[31]), .B1 (nx497), .B2 (b[30])
           ) ;
    IV1N0 ix496 (.X (nx495), .A (a[31])) ;
    IV1N0 ix498 (.X (nx497), .A (a[30])) ;
    IV1N0 ix500 (.X (nx499), .A (a[29])) ;
    OAI3N0 ix504 (.X (nx503), .A1 (nx491), .A2 (a[31]), .B1 (a[30]), .B2 (nx505)
           ) ;
    IV1N0 ix506 (.X (nx505), .A (b[30])) ;
    IV1N0 ix508 (.X (nx507), .A (b[28])) ;
    AO3I0 ix510 (.X (nx509), .A1 (nx501), .A2 (nx499), .A3 (b[29]), .B (nx28)) ;
    IV1N0 ix512 (.X (nx511), .A (a[27])) ;
    AO3I0 ix514 (.X (nx513), .A1 (nx509), .A2 (a[28]), .A3 (nx507), .B (nx48)) ;
    IV1N0 ix516 (.X (nx515), .A (b[26])) ;
    AO3I0 ix518 (.X (nx517), .A1 (nx513), .A2 (nx511), .A3 (b[27]), .B (nx58)) ;
    IV1N0 ix520 (.X (nx519), .A (a[25])) ;
    AO3I0 ix522 (.X (nx521), .A1 (nx517), .A2 (a[26]), .A3 (nx515), .B (nx88)) ;
    IV1N0 ix524 (.X (nx523), .A (b[24])) ;
    AO3I0 ix526 (.X (nx525), .A1 (nx521), .A2 (nx519), .A3 (b[25]), .B (nx98)) ;
    IV1N0 ix528 (.X (nx527), .A (a[23])) ;
    AO3I0 ix530 (.X (nx529), .A1 (nx525), .A2 (a[24]), .A3 (nx523), .B (nx128)
          ) ;
    IV1N0 ix532 (.X (nx531), .A (b[22])) ;
    AO3I0 ix534 (.X (nx533), .A1 (nx529), .A2 (nx527), .A3 (b[23]), .B (nx138)
          ) ;
    IV1N0 ix536 (.X (nx535), .A (a[21])) ;
    AO3I0 ix538 (.X (nx537), .A1 (nx533), .A2 (a[22]), .A3 (nx531), .B (nx168)
          ) ;
    IV1N0 ix540 (.X (nx539), .A (b[20])) ;
    AO3I0 ix542 (.X (nx541), .A1 (nx537), .A2 (nx535), .A3 (b[21]), .B (nx178)
          ) ;
    IV1N0 ix544 (.X (nx543), .A (a[19])) ;
    AO3I0 ix546 (.X (nx545), .A1 (nx541), .A2 (a[20]), .A3 (nx539), .B (nx208)
          ) ;
    IV1N0 ix548 (.X (nx547), .A (b[18])) ;
    AO3I0 ix550 (.X (nx549), .A1 (nx545), .A2 (nx543), .A3 (b[19]), .B (nx218)
          ) ;
    IV1N0 ix552 (.X (nx551), .A (a[17])) ;
    AO3I0 ix554 (.X (nx553), .A1 (nx549), .A2 (a[18]), .A3 (nx547), .B (nx248)
          ) ;
    IV1N0 ix556 (.X (nx555), .A (b[16])) ;
    AO3I0 ix558 (.X (nx557), .A1 (nx553), .A2 (nx551), .A3 (b[17]), .B (nx258)
          ) ;
    IV1N0 ix560 (.X (nx559), .A (a[15])) ;
    AO3I0 ix562 (.X (nx561), .A1 (nx557), .A2 (a[16]), .A3 (nx555), .B (nx288)
          ) ;
    IV1N0 ix564 (.X (nx563), .A (b[14])) ;
    AO3I0 ix566 (.X (nx565), .A1 (nx561), .A2 (nx559), .A3 (b[15]), .B (nx298)
          ) ;
    IV1N0 ix568 (.X (nx567), .A (a[13])) ;
    AO3I0 ix570 (.X (nx569), .A1 (nx565), .A2 (a[14]), .A3 (nx563), .B (nx328)
          ) ;
    IV1N0 ix572 (.X (nx571), .A (b[12])) ;
    AO3I0 ix574 (.X (nx573), .A1 (nx569), .A2 (nx567), .A3 (b[13]), .B (nx338)
          ) ;
    IV1N0 ix576 (.X (nx575), .A (a[11])) ;
    AO3I0 ix578 (.X (nx577), .A1 (nx573), .A2 (a[12]), .A3 (nx571), .B (nx368)
          ) ;
    IV1N0 ix580 (.X (nx579), .A (b[10])) ;
    AO3I0 ix582 (.X (nx581), .A1 (nx577), .A2 (nx575), .A3 (b[11]), .B (nx378)
          ) ;
    IV1N0 ix584 (.X (nx583), .A (a[9])) ;
    AO3I0 ix586 (.X (nx585), .A1 (nx581), .A2 (a[10]), .A3 (nx579), .B (nx408)
          ) ;
    IV1N0 ix588 (.X (nx587), .A (b[8])) ;
    AO3I0 ix590 (.X (nx589), .A1 (nx585), .A2 (nx583), .A3 (b[9]), .B (nx418)) ;
    IV1N0 ix592 (.X (nx591), .A (a[7])) ;
    AO3I0 ix594 (.X (nx593), .A1 (nx589), .A2 (a[8]), .A3 (nx587), .B (nx448)) ;
    IV1N0 ix596 (.X (nx595), .A (b[6])) ;
    AO3I0 ix598 (.X (nx597), .A1 (nx593), .A2 (nx591), .A3 (b[7]), .B (nx458)) ;
    IV1N0 ix600 (.X (nx599), .A (a[5])) ;
    AO3I0 ix602 (.X (nx601), .A1 (nx597), .A2 (a[6]), .A3 (nx595), .B (nx488)) ;
    IV1N0 ix604 (.X (nx603), .A (b[4])) ;
    AO3I0 ix606 (.X (nx605), .A1 (nx601), .A2 (nx599), .A3 (b[5]), .B (nx498)) ;
    IV1N0 ix608 (.X (nx607), .A (a[3])) ;
    AO3I0 ix610 (.X (nx609), .A1 (nx605), .A2 (a[4]), .A3 (nx603), .B (nx528)) ;
    IV1N0 ix612 (.X (nx611), .A (b[2])) ;
    AO3I0 ix614 (.X (nx613), .A1 (nx609), .A2 (nx607), .A3 (b[3]), .B (nx538)) ;
    IV1N0 ix616 (.X (nx615), .A (a[1])) ;
    AO3I0 ix618 (.X (nx617), .A1 (nx613), .A2 (a[2]), .A3 (nx611), .B (nx568)) ;
    IV1N0 ix620 (.X (nx619), .A (b[0])) ;
    AO3I0 ix622 (.X (nx621), .A1 (nx617), .A2 (nx615), .A3 (b[1]), .B (nx578)) ;
    OAI3R0 ix629 (.X (g), .A1 (nx598), .A2 (nx774), .A3 (b[0]), .B (nx776)) ;
    IV1N0 ix775 (.X (nx774), .A (a[0])) ;
    IV1N0 ix777 (.X (nx776), .A (nx608)) ;
    IV1N0 ix599 (.X (nx598), .A (nx621)) ;
    OA1R0 ix15 (.X (nx501), .A1 (nx495), .A2 (b[31]), .B (nx503)) ;
endmodule


module OA1R0 ( X, A1, A2, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input B ;

    wire nx0, nx2;



    and (nx0, A2, B) ;
    and (nx2, A1, B) ;
    or (X, nx0, nx2) ;
endmodule


module AO3I0 ( X, A1, A2, A3, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input A3 ;
    input B ;

    wire NOT_A3, NOT_B, nx4, NOT_A2, nx8, nx10, NOT_A1, nx14;



    assign NOT_A3 = ~A3 ;
    assign NOT_B = ~B ;
    and (nx4, NOT_A3, NOT_B) ;
    assign NOT_A2 = ~A2 ;
    and (nx8, NOT_A2, NOT_B) ;
    or (nx10, nx4, nx8) ;
    assign NOT_A1 = ~A1 ;
    and (nx14, NOT_A1, NOT_B) ;
    or (X, nx10, nx14) ;
endmodule


module OAI3N0 ( X, A1, A2, B1, B2 ) ;

    output X ;
    input A1 ;
    input A2 ;
    input B1 ;
    input B2 ;

    wire NOT_A1, NOT_A2, nx4, NOT_B2, nx8, NOT_B1;



    assign NOT_A1 = ~A1 ;
    assign NOT_A2 = ~A2 ;
    and (nx4, NOT_A1, NOT_A2) ;
    assign NOT_B2 = ~B2 ;
    or (nx8, nx4, NOT_B2) ;
    assign NOT_B1 = ~B1 ;
    or (X, nx8, NOT_B1) ;
endmodule


module IV1N0 ( X, A ) ;

    output X ;
    input A ;




    assign X = ~A ;
endmodule


module OAI1A0 ( X, A1, A2, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input B ;

    wire NOT_A1, NOT_A2, nx4, NOT_B;



    assign NOT_A1 = ~A1 ;
    assign NOT_A2 = ~A2 ;
    and (nx4, NOT_A1, NOT_A2) ;
    assign NOT_B = ~B ;
    or (X, nx4, NOT_B) ;
endmodule


module OAI3R0 ( X, A1, A2, A3, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input A3 ;
    input B ;

    wire NOT_A1, NOT_A2, nx4, NOT_A3, nx8, NOT_B;



    assign NOT_A1 = ~A1 ;
    assign NOT_A2 = ~A2 ;
    and (nx4, NOT_A1, NOT_A2) ;
    assign NOT_A3 = ~A3 ;
    and (nx8, nx4, NOT_A3) ;
    assign NOT_B = ~B ;
    or (X, nx8, NOT_B) ;
endmodule


module OAI3R1 ( X, A1, A2, A3, B ) ;

    output X ;
    input A1 ;
    input A2 ;
    input A3 ;
    input B ;

    wire NOT_A1, NOT_A2, nx4, NOT_A3, nx8, NOT_B;



    assign NOT_A1 = ~A1 ;
    assign NOT_A2 = ~A2 ;
    and (nx4, NOT_A1, NOT_A2) ;
    assign NOT_A3 = ~A3 ;
    and (nx8, nx4, NOT_A3) ;
    assign NOT_B = ~B ;
    or (X, nx8, NOT_B) ;
endmodule

