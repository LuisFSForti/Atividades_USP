* C:\Users\Luis\Documents\Escola\Atividades_USP\Circuitos\Ex1.sch

* Schematics Version 9.1 - Web Update 1
* Fri Apr 26 18:36:40 2024



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Ex1.net"
.INC "Ex1.als"


.probe


.END
